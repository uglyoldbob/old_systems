--
--Written by GowinSynthesis
--Tool Version "V1.9.9.03 Education"
--Mon Dec  2 08:33:24 2024

--Source file index table:
--file0 "\/home/thomas/gowin/IDE/ipcore/SDRC_HS/data/SDRAM_Controller_HS_Top.v"
--file1 "\/home/thomas/gowin/IDE/ipcore/SDRC_HS/data/sdrc_hs_top.vp"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
iMy5HM06y/T1O9CC88s5fTkuBcTGuBDO96rK0dhqiIKavFKxaV8omOG2QcUH0qfPxkvUaw9I8qJJ
1ys1zP/b2bBWwqnxjxPauI+41V9MYtnwI7cQS1kMIytC9Mp66/zUZUtPfs8LszHsoJGdbkwGV7Tr
KfSc+HD+MM/bLfTmsx/YGLblXMACWNL7AppKiFFUWd3EYProJqo6KHYmIHzZnPiIk6Y3LhjYlaMs
A/YFYHmTWyrlOTcg1GaF9XiYzUu3cR4PniNgvJvgVhxIZtdVggeAvXachJAaeqY62+IaYP8O/dQH
s9/kVDaHy/JEbx0s/dogZht45SMsMMMClVk6zw==

`protect encoding=(enctype="base64", line_length=76, bytes=87840)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
yY1QgJY7xph3RHH8nC5O5MDBzobgi3LabRtVZSzf9gRxA2+xrd8hPP1HpCUEaMMllQmKBvKPXJXw
detOE1owVNiYRIRy6KgN2ZAO8z6QkUSX2JvZqX27DfhIaGdpZQ3Pw694cy+4GY994r41KNTXe1hD
MkURauZzdfy2etwZ+eRmi4D2No5ht7naFvPpb7bGzFfhEoVBBp2pSKaA21IiJb/WLO3LLhOJl0P6
F8G+vwppUf2U7oSrTsTWo2ZCus+oT9UufcYfHY6M85mDgEcLQUj2b4e272e4fsloiIt/e+3+DqT/
sl/MX3OAUpfTnxUut1RHU2Krnyf1ubHfQ2VdPLmciVFR99K2WjZNVKCs1BxFG336Uf1p1eMYLkeX
FzEogCIyRRTBVo+B35O3ly4Qfllx1DVSnDD0kXesAWJ0qQgagreJiLPlg/MsRM9hlG8PENwws6qJ
FshUjNCMzmucmR7UcmfOa6zPeMLGjVmA2GG5/erXZGMRIyvoZqIeVpdSVLShE0kzB3WPahcGb9cX
eXejOJLsjJitvKn+VBG3ruDNzQOC3Om2DeWGpIB6J7hWT/hnvQr1X1MQdCn/GU2hTzgIowWzqVMu
lgGn8CbL65XIE2fkRphlyNsttcZX/qs6ux7OsMdcd+5LxrTYx7OwYjciGVSRIXipLhQnSDADBqLs
yYup+NOhEVQwwrU7W4CZCVZPp3UXAZPwMBmSQvvRUuwa59nl0gENcx31o4p+An/2wu1FOPf5an6D
kvi8qKGKWgbHBr4LDtxK6FwJyYeue2oDbcnyOY1JRRYNRIq1wQio/sLOuMtnpQSa7s17oHsbkK2P
gUABcgdalCUs6gV3c8XjvZ/h5kvGV10m5cYwehwoBWXwtf9OBqFfcLP04YwDd5/M1yUIdEVuvFA2
Myi4HM4gEdBuzkRuKusmsMxdUQl8dlb1BmIbyTQaxO322vGxcv3gZYYdGAykorf7mnkhXRdRHLyS
/LjTTce5diFG1PRQZzdEUjQksr0+nqTn6l4GeKLtwygEtSDMwy/Rtyv9IfSR0QP9xIeIzk/SY1wW
MAPGcnFp+Di30qGUOo8UTA1FmTR3N5A5Paj1tpCKu7+S+9hFkGdes1RwlHerajZpHVQwTj8AxVWp
WSYk7Mt3oLwMGn18tdH3Fsvb3AweWQlk/AlDw98JnO5ZxjjvD1thckvOs1KlmluhWkEq08oKCOup
7caNbzPDJrEldE9p5ZAMwGPBp6BWBszk4nlUAQ8d/+e5VyrMK7la8TtzWWEC4E6X/E+j4Zv6+2/y
uyItxJhAjQr3G3Z3d2eRA0W8Mi44bAFfraobmB12nRj0OexOdpduqbxHEFJVAo59QIc8TTIbZzB0
Ge3APsFkPqe9RC3tnRxdM6HS5TCtboS5x6uVxavyLahlmjVttF8p59oDdc/srh/jIj+/8MLD6mvi
GbfopmQSq8s/8mdQ8c/LITtuCOr0zDgfqxXBFsWpi09WbBTgEKl5bT/D9qC+uQwqFJdNks7gzTCN
463LS2h1S/znD8nYRf1TYA6EntBsVrGd4AejAXiC9BTu8NHksnbTRF+JuUqno21V1E6XGs23kKGm
AxQlN+F4IBjTpAPlUd4YIICMN17c1c+dr+qt4sPhMLpjoz5v7XNz/URAmoC+ZySJY5C0VQdQlVMO
UPqA+0sNKGGDX17VKbcuRjwIRu4RjWVo1NxgwicMq+V2uRzqTszkP4v/FnZWXl1o49Y7CB5atpsU
eCq1Rnrrf+tbs/QfRrtH7D9klsaa8/wse2ZLdudvCzrBEpccSP9AXVpywI58iPc8wEtPcotza0rX
WY+jRf9MsXwQFPhF/biSH4w/r9trXfMyERlwb7n6q1Uu0SE7YnpwxBamUJXucsHTQ1xIJXn7euSP
E018rPlY7lnK7JoOZ2nZmvVTyDZgxr/9AFC/E4bXHkQlTdAMg70lbxYUp4lQMslAGGix6DCs+hFu
+mNHLmr9IGOw8Yptb52dGqtEdMp7l7yyrLImrSu1QJo/qWw0+T+qSp+XCQdVXI5WK2qaxQsIBYOS
JWyEkxB5x6an6qWLvwTL8N9YLm5m+tApHHLOQkLT3SUKFwpU8y6prtmDX7Ac2TXwXokBSLYy5IDB
DRD8oSrmIi9GLZZ7P3wvElWfb0jFEKa5u3TpOhydscdO7WzNZIISCqKzwoj/yrCz4xmLT6FdZlj0
UWKLFn1Na1bsiUGQiDOIEXT8E/rHbrrvc6gOtJrUgO8i8Ydzp8645CQCeNDO7O1rVGRllTxZ5cPe
VnTUhLyYiT7LUd7JydxO4MsEjFQLqUhYYpDHbCWL7CpoEtzy8Ip38yLy/kR2l+ypAUh8c4gccoHe
Sh2kbgZLXDrCB62AFB17bUm4K5GKHSt/7o2LzvDkD0wvw73TMEhhjGpnCmnMysAlMtniI0MWd9wr
o5Fo/0MS+U/GxQX94jVGWNYPIjo0BQuh6E1SjVLqPUBzAbNfSpu5ixuI3g7DZBe7w11nxDs6mJuB
8bpYUn8BfSPEVc6vpK/FDpwVCeAl/zQcH7Tcd/FuksG5lrcb/RvNi4cV81bnJxbgY6sclbIVVmF8
d6WLB7B9kbiDre2eQnq5VLzz61lgBTwdC9h3MNV9CvIIHvEtwU7fZ9ok8OncgYX6GVN8UtMRt5H+
jkh02WOQ5ASirMQSVvQLbgd8re0XEouEjbAPFWFjE34paUDw6+XMh/NkOsCTd+MDvynI3zpGQa/2
gbfw6w76NZ9Hm+idMvuuephp9UzZylGdHgidIccJjWb898VSGsku6HtxFF3G1tq62i8xGbYev409
PQ6Eyrf3Vff6Ts4gNF4M4gC7/hqrDCVaHxoV1YRDdDfEdysUbyPkfvBVkOAC4yogjjjbkmQqMJaQ
5SV2wFiBN0HLpbYd2Va2ZYv6FSHYkcnkA2jlZ3li8ZE73k5K0PmJTSqJk2pENGrphZdUgTpER4p9
ZQD73OJ+yUNZz/HcUBr9XtnQeh5M+m0ahrAaXZPbszTiAY44/rXDYK14Ww0mUZYL5gsgTRfiBza0
GvMC6TufGscnYK8L3s9oEPDRSz/p4h3xm/DoFAuic7tWK55IsuvSRf6rdhVZfBlKKdCLPezecQZY
qjGpsvPkxoLrDhxa0ymg4OYFuUGKtOGwmDnmf4bfXBAuMVvAGYCTLImzwzWBOQiJmVtmD4XJ61gq
+GTgKOnjOWuWmR3+I8jZvimxfbSj+fingch2PDCbq6tlTOMq6+Uow5qO7Cs3eTzh6tJT5BBbKlou
cUdMDr5Sowxaf881Upu49vkXbC1VeoqoUHoXZGq4bqkLwSOrDjSKPl3LKwU4LFSj0+KW6m6i6dJI
fFNUSwmYb+K5ym5tH3XJysKy8FT/UEg01QUcoMAcJpyHKcsf7z2VBJrD75yyqyYEyXykXWTqWKvN
hw0oB8QjOYf7MTAyMc190XeCqcEGwDhVKFgcI6k0NBsiEmH00ArrpTKVkmBkupM2wsDtyhOQ+2tC
Vxgx4eWISW+iwfwycOPIzwckemfekL4nXvOh/lAutBNXo6JkFPFAKxq0rYTl7POZ+D3HsNZ8m660
NQr5X2QP4KnMiStHKDCQ8+uB1yfxGEN1YOV1r+LqfMvKlX76ZEcJijYco/29tKruBIQBbWt9crC4
PTUzsjxW98fX/UrBZAcExJ2+Gq34If5ths5wGMb+NjafPT4Dm8wcUs0SXiHgb9ASHIrpqgO2mrQV
SkafzHJFMNbfpQroa2E9+WdPHGrq4R1vs+lE9PLiDqZaNrqaRCUPi/1n9qJFMWRc4AocrPVQVK+O
qpxWeH5ppAkBWAmEvGkuU13raGzBgZGHVsbVY59jxeCHkQ7FoZihInrIoacIjOuS7pRzFBBR82iU
KXYgWtbtxDzHQhGOJXVMMlnWXP9EsdnqbFa6DU5Evh+/eidfyiKsphYd0wUAPUJXK4JTHwEooRb9
sV2/B7gpYBOdVcf6QXRL9PcstYR12rLgEwS6TPZrVq/J07cEmblmDCGcwwqSvsFj9qmr/vEnn4Dx
a83xgoq3NRC9vqF7vuf5J9Dq7jeZePwlhkLzMvBHKPxbVa3ClsLkZ9iV6Tc6N2rIQ42oZRJk5bIj
FHXIDqYOnGxiS8LJCfQdc4sJfVH+6NHiGMeYat5SLURWveqAXEpnLReHyxI9yvrFFyXp1S/2aQWl
dDkeekCu2bk6OLOUn6Np1DBr6Bo2xg0ow3pRPwjJv0zJRvAbls/43VRhSDyN6nw4rWsjipiaXrv0
5HvVHwiqHr7/smRjqy4P0yF15iquq6QCF5Qc4ui2O303e3QwJjo2qH3FRE3Ya6FfSPWDlHyqGSRy
JtMXM7N0k46YZ8Xxzs3iSP7Bc8U8f8x307fTrzn1JQFpyeZilF2LKi8SH0kamR/qpPnEPLaGly6m
0Wa3tboCS9uM0N4fCpo5ixgAOJF+pT/8a6HwHfma5/Autgqbsr+tQEcearBjiwMRzUwsCpACATqW
DfyByoMAt+nFfKuQdroV42Riz3LhiOL+T+ve8Vc5dm50m2GsLgx3Pcgx1oIrPXAXimwlaNg/h7df
uu0CVEbils8lPBEUI+YrXzbOi2XG9zYbwU8i29CCodREPmRXs+KnWOb3v77CNxmnaqCGnTIwdcCW
i+Lpq8tzW3qKFRGM/szh/F85mCa+fzEtfQzscu81CV+SONBj5yzxV6F4di09Z1bYsbyNS4lA/hrZ
fP2cpitF8Yp+yEvT1jmwxgVVjWE4+KhBZp/j3h8HEc9QaZS3+1fmGu4OZfTsYNGrzeFz/grOFbkn
q9I/9TgduEA2kf+WhaUBeXf0lAjRjZUu0m26iysRRiYoeFBZ3NgEfA1Bh5S3Vs3n2m7vHCQ2afif
J9WkAZROrmF45W42cMKoUM/gPIHyDDGSLc611KbDPaFWxH85/auB9mhes6zhURGPh2Qk3gn3TeNg
RUvTfeVZ9st05m4cSkrolyxesc1I9rEExn3Y3Xz9eVNAuseYDOfEf3FUVBMfzzF8Qkf2oLjEDKyg
JEp/FPFr0wws22ZM0Roi0IVCXKtQleOi8PcZyIir0iQpVJf3cNjALRBQGoBZLAUDBuYTp5XmTnO/
dNLaupHQvC56d6wJgnRlb88BrxxvQdl4KGg753qVg3nI9eyt/9klUBCT5Dxo2vp7Rl6rM1EeTfTL
HX2NiwtREYPOc3m/ZfbMSmDyf8nD0a9RDMMsPLg05F3keYhIBeD61a6vy2z9hQtYoaUgWMSC3x86
RWiDFHsLVrISUtkwWdqmsHufHseA2F3oFRucyA4+VQPAQiUjX+iGEBJfoStfYXW/xzLNUsMVEseC
ygnWVKrZTXfg/wuYzGvL2LUoixWZI2nl5oIRYT/WGkSkO8Xa3DuX3oSD3wSeF+J8p1ZquR8HUWqa
07hkcu9LM4rXtvZvmFqQOtGMSauBw7IEFxsqxm+grtSxlco3Im3945DvPKZR9WKp/fawU7CwYAKF
jVphul+YFPIuQYp8m/GeTcynJUJAkZ3R2WSw0SY4KsfAsbIRHzVXMJl1D7bDydtUCN5A0WxkUF6H
faz9OD+Gw64ICKVUvCOwdo5WXJD+B3wvmNx48qLtQkgn2NjJZrMjYdUE7coA2tsW1tF/TKSizYU1
TTfLhDyfH60DQFBVZVQhIWFzKv5nI9Ayc8ddzJhD+pi4fncFrKtv9QT2UHzIaym+2a+wgSaHPT09
guz4dBixErzoYw5fZJvaSjlgh/fArUo6Rt/g81cRRlbmFyO3LtQx9GC2v44sFXWFKaiV4ap8sri0
eRo4uaLiEtKx86hhwrmOvn1aPTNDzGefT/1W9ZsKYblrlD96Q8uw9dQoHcKHLDjkxFl1Ac8pakqj
P2hMgbHfqQAmUhTDsya6gwKbJrmmExui7rRDHNkrAJ1KysBxDiYQh88NM4Bpaqjsbs/nheyzjBJe
TgqQay+3r9O2X7eqhZDe8iUcf8lhvrJk9Xmve6YAAF2ateu+IvNp3mi+doSRmt5alPADRO58LJR/
IxLztiN8DCQQe0W2qFgumlkAgDS5iHlrWmH+1jnFlEX0C7FNjrVD31fK8Yh3k2a43diBzgDrW5DH
mJU5Z67vhDqogrBXmJgknMI2rGziD+7L7ibT+TieEIbebXtTj86mfzQPNlbeevWFHI14hRRsSNmq
Xa5QqyFHDwTJ+1/839HeDVfJyA7OVa7l1FSkPLg/SooIU4TE5EfrCaL4jAnDKdSOO5c0Zjy74H7q
GKIopMO6HpoRdSghx/fLfQ7WrkLra8uULRfFwr2E8bCipMWGrZ4Uvewa6kYB7cl3TpkNwr//Nocu
0hCh7LmNNoFP+DH0ElMJSdVLaxSQ3Zr/YNFpQlcHwaKmAGz7NqiOmoQJrTwCHA0wELKLW2Fqc/8m
fxhuBmOVA2KrbiPerSp/rSakDD6MJrJtrFiqkKQRn/Gpw1hvYTU14KXPkoy8Msj0agJd8l/ekSFS
IlhXA8ZM0YR39FodS1rntlAw9SlC7LBfmqMolBoRnM6+C+m9fyOmrEG2gY37Fuen7xtPBrcQcPVP
o35dC19KUMWSxd4swFtTYk9oepJDHQYP0hw+prJCrXvG7cU+XmrMw/xulnO5KT1K8/arM7tG1DFn
sf7dl1IERKDrKIPUnLCG66ZsC9A8M3XtviM2PEI0j+AyLQxzouh5PoMp9DMSmnoExco+KQG2Ygx4
YKba7ulTCEyN4BJprNSoHCnKobYWi6iIVHsnnbfpUjuFYHAYyfjZdnr5nrp2gnqxHacvFmJKj2jp
cf7fUkI4Tx3i/ydyjlLFdbJtzfjRhfXcHthuKZQxRjAtjvQc2iNDQogtfi1ZbxgrZqcEkN2r8MQQ
YIv7X4viPrjouXNmswUYwcrFYv95Dv8OGhnUi2BDW5rpjhhd3U6Y9EcztrLDDsSqrz4W4qlRgID2
q3tfEXl8yPvRRnoCbTX7ShBiyenHSbs4DFEiLFBHlmZYrMRzMr43l4KI/d4+Z9yDhMNbsfIRSqyl
hY5Pv4aVzj5x+Gw6YXHGyKJ2etKEQ3ZhoFXX6dXGzUvs+2YO6beXD2z6E1mM+FEQZlNX4sJSPvCi
zMUrZLxylIXMrHJ4Ems2NpmbNJjsZiTrcshgloNCAx50VGpfCktFGEaiSmh20nIegZDn24yBu7nM
39jfpySCXo7C+cnZe/hv3WjM19i5oAWyYUt3VPSmGnDQU8DCv54uc9od3TaKRkHb+A0M5scicjlM
N26RD23uLGwNBmSs9xgBpymwitik1vosyJXDQVxMaY1g1OafnPQQ94Ms0snAFFpemudzyi3YGlZ7
QqZquZpdQmZUUsv/G8KA4Wpyq5nSgGpLOxTd9MQ2uTX+5T3J9r40D12vdjuiw/pXHzavQr2Nq/R0
SaCeLcu6PJcw2Qut3GjTEcJ2QBRT7Dhtbp1GP6KRqj2VMnbU1r6RB2+oQDAw/vWNn+Pcivyf/+3z
B4rqPDTGmHxOuY4QevGq6WmsvqGgNZuWK+XqrcAGZtZ7+uPrFYaXcTTFp6l45wU/wY5Jwit7eOLJ
V4c3YUZKmYzr54elAcKgp1QiEymINJK3R+XaIc9alQlJ5mWMYNMXd6Y0GTARkTQnF2w/NgMuF2zh
uQOg50zu1coU4qkzdJid4g2dwJ3zRSyXEqyS6cdglsFOR0ixtd1pPdTZOyd2X/9SW5E3My00gSkB
B4/j88FV4Y5aQ4kXwwBX889f2/0rXcHo9l01hn88mcPTKH2CG5Qd8nJVR3seoTNFEY45nwOH3Zmn
PnVwHhVEl6RTfV3o/SHbf2l+N3gevsOScdoiAl9ZNEaZyPd1KTO4q4FFNev7xkLJ+yYMzV6anHci
pgbcS8ESSAp3AX1ZbmS0JQXK5r4bQyd81yXk45jDXD446azty3cfLLWiFhaix1DS/H7IEGiPa3Au
3FIFqfJ7kQnwYqkopDPKtdLyaXIWSn/zVr6ttj7haOj9/WElpNbbIRBHPzc9Cdmf59wKcwnUBk8x
1ILCe026nV41txxFiWdXvQrVZ8SunUIm1Dy2UOku4f0B3ClU8ZKnc/4JXYt/OWlbxexk+S4bX0zC
Cl73QhgtUgl5tdHcTb68vVTp3vZrJ6OQa69ef8X7+lu/M+fT/R+GIzUuN7IDA+9KtycK+SBqRNnu
NYb1zHgCcoT0gih4LZre9GbKYLEMKA8xlBIO/vQkYbejLno1b04qhx6h+aZD2s9g1zkdCEgpdrKE
q64VQ3GIcNe61l/NauA3uCWZAnwLMw7Lan376ZpErpamUB6TlA8OYdGc17+IkH3iRg9eQP4TmDQd
i/AApmiUk76ew/ugBNMtVl1cjYgNrAtdXAw3cE+DKwn1M/5d0QI1rMH78nczFQ8AtQ4QQ+9Pnfz+
WihNwL+ZLBDrEEF7Y1eSKNG9/MCNOhm/ITTOit0vdWdOekdkevTbizfd9pvOox3mz3GGzQ//rksy
cxYNAR9FV/guKfxjrUXbxKIJC4UaIMNhKuQ9aIlUgtjAUny+nsypbvqYIx+EDNvGU1sXbM3lgx90
gN/fb3pvCMa55ujNzoefUZ7nR+fMEjqEwVTuKAKW6XcHo7rmmBoe0rXtfh2l0fbX92c143FAtKIB
ao6VIIoe5l3LkdfnUEtdsrFMq7HUkx7mzVRfLrc4BTfK/Qq2QIIJPqhks1PXFJx6eoK9fi5gzEuf
AG5IRju9A5YwcJpQ5USY9EjWBqRzIgy2RSJPsD9qLIzGpjc3wc++CUEGfE7uwnck3O1ugjYHaMvu
Se3R4MvNI/VLFmTe3iMjRO/N/2OjSYtInhIi2FTYVUWNdYH9JESir7sEKWCnjApfNClNGuzGOwNb
QQ+SqpLEvbzizS4LbDUQBiZwCub0ZigrgrdpDTwtkNDXBCpThBRfjWpKYxrGrFzJHcSeQw8r68Db
AJoNpzNmEInAvd3+aqLBCOGnRA1G4Z4x1XFkeh3HZOsQXKCfl3kGyCsXW8p/KmDiWhD+t9ZTPejV
CBEI3oxcflkT5YY8BMYOK19T1bvjkBccQabgXFM7Fs/VBU/hHPjB2Rb2HigJOh6hsiitVLckIk7A
RCpVnm+qOYVewTXOSHB81A5xBSjv6Sc4j7kozkMWTLyGp9422CZUy+VcVPJhex9YG6sx8tYn8WYl
7yvniqKP2UPmO/3GuFR8a7KUerG3h55cEwMGVZ8upXz+oGJOfmD4DqYR7b94XK0OeADC8OQGQwyR
/tuir12Qp48A/VljzYXCGmiwRs+6jlgQxprtAFHOA5TY5j3Jb5026ScKy0mHVCzhNQcbV3/4mU7g
i0llo4zyefLWd3dKRTmmldDAHjj9kBCToeBXuwLFILdN6/dy89SIB86xqwjBO//h8YpxIqdYYAmk
AiW5Rq5axNCIn2DFlK36EjW1v8zRoU9+p6ueBAH3EbjoSOMurM54dk/tG3Iow1QFmZ/f1GJMCrrK
LWp30I54w3GeRTAiOkVDr+Fa1oLa/vnAs/0uCQGwAJm5Ix7f0ntcccBLOsEQO+xoDea/tobtOt75
IxaqQk806kLrylMF50ts6QHW8O3i2dveLb/TVIindn7pSbp3mYJwgrxQhP69meYiia1WMw8dwDuU
uewy5lypOYb5n682kuVzBKcnEOz7cQapK3pwhOR5drEhlqFGlKarxEy3KO3wrTs3PMVZbHHkxpvG
UAzc6ziUQrBA+i/7cDOlgc8xQ3aehc0HNMe/8uEmRc4nkc3vlbDSQ6RsutBaPjjCNc4jaKw1CRtp
HygrPX+7C8ibG/BeZHfyvSqfWpjZ1kfa27JC2QxDkg6RgZB3vfasmSLaqpxCpZRa0HBwki2zZ02l
Z6F1Fiji6T7gLE/pz7dWdUgw+JD9Xsvq42fs4wawxajHMPuSeJdYc1vzAMRH6Vvxr0wJsgRXhQAi
z9LZXpIDS8ibhv9wbQdq1iPGdxZv1nh9W7EscliBypc2n9ADpsGKA8UF1fL8+yJHr1qYeWrZa02/
hQKTlcqnqCWdBS9cNcCsgeJbiqlzvX0uLCD+WxXzD2MPHi1C1ztE5a6yfG2vot8EJB4+uVrhDhlE
G/xWGaY+z6OSn66lSYCv2Uzkub9K5tB18Bxbc53SipfjOWsDg7DXJJnUfKR9Ob/6D8OlRF3N7ORi
NItXel1pHnxn7/G1NOrB/2dHJfsktzd2ivqnMIalgH3qlXEeENA27vob5RCju0l3fMNBfgrJK/Lc
nqiuVx+yL60T3Oan/pqNiCBI+T70W4jQ/GF8AqJkpxSf5BL6kJGD03OUGUO7Anb7gzdaBu0Wpmeg
R9Mu0ltD/d3/wmEuNMxM/OeE+WhY/gQjfsCYqjcSXp76Pgd8abvAXZftY4nBGcPkXDBoU3BSmmly
Yaa6e3vECJRU0c5DpMLqZKwmWSsoNzOSmzW1wklhIaiEbFhnbE/CskjP9Szl7RMOU0xipuB41EeQ
Vohniv//qjsfrkuEx+ym7ZbqwHOFfY1Y1xchekNQ0zr5a/x1KqmXzZhmN3M6N3uaLuaSrW9hXoAH
2dYl5vmbGG1VsMwJvRpbBLbYVPFrnpcZwWRWX7dvKWHgZXUtYe77WX9mGqcT6qAP4brbdvhT6Rqa
J6X+l8RMCGKhVD/jL86V4whyhpI6WXv7V4/1GLid4nfGNxPe9pLU6T+RtnQDOAjxoOBNUflS0IeT
/nb1aiMXnQMOC36ERqrjGiywCKOh0k7LlnvKQlPrf1qmJVrr15sNeuhSzPTIDpJggT79NpGnibMA
lkYl2wqVvshWixz9OBCc7WLe807ZFdhhR3sPm/ZCt0X+WX+j38DIp6K4VnQoTh41pf6tAT1ZE/dx
VDrFnU4Rt03JcVmfMuFyYxua2ANVL1es9Bjzi2O/YmD/36spWTN8QThE+FU0VCERLQZBmeVxZQh/
B8zv2ntqxo8x0OwlLB1YbMvk6HKTqOpyexG7t+Y+0eqbeECP9zKKw0mxZYnOGMOH3bqDkkBuKBWf
bUPADVIl27wXnB79vDKtx/GHaD2L9Jrf6V1+3Du5v7zvaykynJ3Sk2RgBq1j1J/snFfmhyFj9Xx+
HRJMA+5MBFYl/mi5qpvTD3AwcWM1o8MF7CQpjcI+guIky6Ympf5LKbeuwYcBz3l2ZlIHZYRUyT9P
cGcJcxN2lfDGoiolm5rEZRt1NOsYEim+UluWCPsgcoW7drgNdpS9Gv/wVXx/kLzPJ6eYLhr6MAIH
a+prehBbNH+GMztVFtA9Tbo2aqxOzDtdT6uwmUcmNRHysEPDfBVreuqDYKYI+eSwFTJXPfEMVsyU
TxBl2aJ8b6lCwi5rFCsRH8d6mGyrJxSN8dguUAxXwaGiENSsV5o/+Q7Snlwtr1Mr0hdu1OQOWtnX
6pHIuGOrWVrE+cGoMzWf5DM5mtBNwlPhx3pvhM2nBHvy//rNrDxVHUV7CBmwxeGg/n5xZzKGZHkJ
54yorT8dXckoVEeUluIlBZbtmdtkII4p8zYmWY6sWI/5+m66dvkiicHm1P8P35ft67eRFbQ3+Y/F
5g1+QxfnWXUu4hebFxYa5RB4/FM7nvrh0bV3/FrvasMX5TWawzdOS7JxJRjezOTLKaYm7cx4dx2p
IZK93I1SVy0Mk9DJzNoSvXqL6q3PeQeM5W1fYhWcwVXdVSO1ZPK16SmIBwMhKyvRzabIF8zNrTve
cLNyXnMUXYmATUoEXvDsNLbvPWT2X2ciUv6kXhpsnLShRMTjtNK+MV3O8LF70QLA/bmNabql7f6e
OGcKSrUlqjEzPkwRTDFkYNj4XfeOZse5xMAQgBJwlPVb8CEDyswKWau5V4X7U0gWE1XcRFDE8tVR
O8ynKFmx35QweBVfRrcxQqNCYkumz197EBxtSKfYvSuqO4F9ZsDdMziWDR3lzRRN/dEdomdcw6us
sDud5wMz+drGlZzun/JVmZjNKpNceBodRJiM9UQiC2UiB5p/RTql50czaQ0PFZnR/3UH0FNWEEPq
epSOi7X61O34dYCR1MYrnxiOPmI4K2YvFE/A1RxkTCPVVW+K+OBjpZSA0kBdEGNlEKi6YgbISwBp
QKPGAv9pCcS2nVqPBC4hNDeqkh1gfVkiQcWq2yO6zfDY7EeobpImmlPNzU7z3R8Jgm2zRXaL1fiv
c6PPkU1Qa5J59AaqlVhZ02FBpe6ViRYVXnQ7Gu+UdogAcTQ90n3KwLjQU3T93Q3LXsStHam/O178
hCpuOhBSNdXMNON4w5u23qfm2l5JA2RCe+KYQDTtiWUBH0e4uQOvz2GpmKp50AA/KXaaWfT3pHjE
Jv11wspu8SNkmq6+a8FswT9GO4WQ3H4IDWIrIRo4eaURp/4j6SReIiOTkFXE0VkaSUhda+4aTgOA
Dv+6/BGpZMjjCo9Gk3YmN3bEy2038HybZcesXP8SgGfwJHI7njigabrSMec9O/0xjHz9upBfhvbm
21Nc/RSPlNkfYJFuhYt2kFiOZFv7/RC2jQAtJgvHsWX7UBiBRGBvO7eWD+fK7adFvK4Oo0Hye0T+
COEr9MGGGpi9Bzc0jRNVX6IZg7rTGCR1WJdcqZ+UVcllHZRd5jVc/o9NqCGq7IcoTvVmN25qSetI
tV9+Di9PDrnGAfAaUulHsFTWTx7k5fPySVLfoxswpyoSxaHwUYa3ArHyKpVvzZM6DTNaEzzO22H/
SPB99fW+zpoDUfGSeq3ieJICL0+k/lYUtPKIBlveG+odxXuDaanK45+mSJZrj0T8oYn7wXb+YKle
59hakeXqDasgEhUcKVmYzbAOdhsXk+1iC29K3tLzD0bdd7/etfx9wXDJYHb6/b9ZY6we1fATR3hV
FVtRT0dpi9Ic57XgLqs/krQSiTltnNnAy2UrjMq4HdAXmsOosz8f8nQmPNBl4hL1333t1HaEucpM
aRzHqFgvY/5Zz6MDuYCiG6GZglgQxh03W3ocnakWNxlrErvvq6P/tkbJpLeydib91NvAgLHeFm/Z
0Fv44nN2r0UifkgCf1EyGy3ZDlkM4fcARyzq3dGuONnctsRlSTx+nvZf5ZMbyiegS1Ih1Ngd0RAV
OYvFGmuSBpXzxYcjdncTjlGysCY1TKRNIbyBhE7/RS1Eei7D6AEh6J7T7rnHnOcapVQxAbQW3Ras
o+IbFLO2aNciHPHHs0joYKreckON04RyDoLcneHmptAmRAKWqOoIr2+cnSp9mmnqNePAokXSwh/V
8n7e53wh7/Os+MTpFpkxcHrlkJUiM6qvYG486cmqMc7Wkz8mdT76OlZAE9IqOLQzNteFiMZPCwcZ
Cl5kuq3lXVYZmIfalB7TawxGzab3s4muZ/IOMV4t1ctG1BQ9LQueQ6pzukdXrlAlBjQnvIoe11uZ
UJdy9Sbn16g1KEjU4lKP1HpdQSLvuHzQ9gznfItXh5VoSuU0hBPLtglQNlSh2evhZdWX/sm0/ToL
flgbub05xEF7Fy84USbVplaJDs9i7YBuaascVgi8G3w7Ot1DHeZ9Oha4TlqrFUdjzSyTpXvkN1pe
IH4lkkj2Xw3PgShjx5WCuxLRQGy+Ma+BwkiMzkQk4xVxOtmq4/Sb/IFp3G5zPf8l4gD3QngjjTKo
6Bym4kkm4EjEQqkvecihLBhhRTQoClol7KSWeiSCUb/6LRqRIJ16Xjzn8LZiSXAsjWAZLFeXGJV9
OfmyHK8NGQUVBard55N6NJMcMqScQFazKjeKV5AzFBBAipZzlBYq5wQoBa9Wt4Tgg1z8uinizmN9
RTp7tUlK0XZooVSCkL10o2L3XCWlMutdc+46njDJ5skMqmh6xUq7NraKaegHN1lxyDCDJca/R4V3
C2ZEdWGTwcLJXbZoqzzEIZf2BSv/2/mUQ9od8+gVi9SIjH1gu38CWgQakdVHQctWfYbwcIndpNPq
Yq/UQ0KeItl2YTqcsgt6D0uLSr2FJFemvI2/nOzg1Hsn1qIGe666dd8tp+3bsddD+aYyz+UVjunr
lAm0M3Pa7J21kkDp/pznzwd00tp1vqeHF8EtQfTNVecjux6FtCuqL2lJgNe5KakmPAUKLC5ej3VY
U8WgHWl7xy16u4xjn9yVO9wB5K+sGqzgDEc63VHgLnN8nIuxHFpL33vtqY5iZTa1X8eqnHUt26Mb
L9DHS8xD1ITSBcHFEl3hm1QiY5V/NolSuLO3AMqs40c4tyfuNswFTgLIlZMl5ETHbg6o8mKuu4E8
MTXMdYigbpCjSWmqMRDh1brOxZrc822SlnyzWwFhWCYei8WyUAoMbEvdSWdmjqGo+rJqxXnyz5zL
fJ8PAZbRrajkcoAoQTY2wq9GFYCHQERIe+O+UtG8he9SbiKkOZMYgkZ0036y+pxvCTEgmmfEUzOj
cGdmNWfgLuFsKHtvK3nuz3hD7xX7wn9iE+iD8Zrdazf9WBRQry2DISWGoshvKWj1RrH6l9ljFzLc
slQrUbobLCzuGq87jhwfNwhnkDJtu8eTT1kcOh1wnVVYYf4N/mNGjH8Jzha0uZrNgN6d9UPRgPW2
n7btxj1uhaE9NET9uTovU6Nv28Vo2wMOx2myn7t5yyqW2ip4KUoqesLlKTFlT1nnveFr24kHSFdB
uWQVSYLjdEQlfpbMHQJUskvNnNA/vg+pqu4fsmyTqMxsGW9P0Hs/6NiIBtTUiXYpkEgu9kj9ITFX
OxwWQY7XauO6iThK5J8pEBT+0rrD2vWkhZCUtqBCcdKmRThFs51Adh1AuS0AuZuJR1zFxrGCugMp
4syvmRIrekY5Zv+ndSFD+RadBT0MY6r0iC18moSrBt0C5aleltwsR5lJO4/LJIjQXimC/jhOUIUX
uWDNgzOb8LmijGh0crnE1n4A9u5ndh5yVK4aIvn0V0PuC+6w/oWP+oRMrO/3puHDtP0STmWzAHSQ
cN2xaR0rxCIN3Mnkv2fNE2TfchjqcpyCEYgbqvCWsbwIJb+6j4bcdEZqUuhzfjEa8EPDeZer2k2n
VV9XoIkd6/DgRtSRTVHQ52DwQmZchI6t1XOrCYd6RMZmfZn1GIgGNs9DT4RVjHpDRENDp+t7pV+V
cJ5S3vTfqwooE24x2CMngLQlvkUlSUUtYnJwgEzrAnMLenjyRRSo7nktvrOB1ngjZLxIrMW1BDdk
3Z6ShXxwe9TCICgIR4vifrZVX73ML8+7GccGlmw9soO5zVp3CUov94cHf9oNtkOrLveOE1TMmHaz
cEFMMouE3HvzbSRBDpfAvZdL8CJdIQJIC4HKsauKK2onKZFE4hi0gil+ELP9dN9aEtytJx11BQgk
kqdOEBoppFlI8wZrhV0aBpiQ1km8Isqm72YbFHwdmrEee+9p1XtaigSTHaX5xai8SAe/5hY6iget
NmiOemP8oe5YcutVuw+PM+bCYTgWgLJUT3mQY633DEoNC5lBku2DuPrt6RO4LqbySXhO+yhRo7zZ
+Syf6WHtHHsQ/6sitmL9r3OyWoFYVM4ZGMZxWSj1EVPnP3SiFktySfVWJ/QCuuZc9/1bY+XTlbA/
m//tR/jMnLe2YsbAmbfwW7zKeAZwhsrsLhfpvisJD+g0KdPg/GQUiRwNEGxaMHMmKNZHDhdUIlrj
yjj5qN35HLlvAPmTSYD1UVMIj8f1H6So9sD9E6a+k8NQydUkukEDmwL1vJWg0V986fZumTL571nK
umqG25NrY4Fpg1zug126EpAheoF0Bl1dA0x9YhWXbZVxJvbNgYvo0o2zA36pR3g73Z4lR5rLSIkC
zkDlhm9STDPmWXMGB2aSOFpTyQMjUoA3Mma0Zx/LXk6tpRNIALEmyDEXZQPdgUaDbMYMHx5W98bd
++0uNle+91jIr+F5arE8qC/gmYVxLBQGMqcExwP4AHmG/nZhEV3Xhw4D1yrVo5OVpCyhEhFwpxJP
M96+DqLrAUjLVSpU+cyQ/kVSrQDrZSneHXuBqrXNYKcmJIocBobzXr/6ZCSicJ90EJfHVzuOoJ/Y
pHMGm5wGZHJH/tLDvBJjtMtjuPcpCVnwWx6paLf0gePk5j/94MQvLEXfZHYSJud1E6OXiQUqacbR
i5FBNBGB3PtBoc6oLS3v622lV8Rz0Wayhdv3kFFrYX7jA6+GJ0wCCI9EI8liQNW0eTe/pJ4bgaeO
VxIcrWzAYf238RfFJHKo7X+nWb6AflapASj2EnWn3SuEvH5XvWHGedfw+qBH2NdXYNl5nwACtSwF
p02mmROjOQrdhmLVAPXLgBlkTNeEm/kOQbdL7xB77PWk0x/yN88dF5iUDPr+uRypjrcLzdrtAe5E
JIpL9ynHl/SdGUqOKhYTvnbzLL8JG4UEy8qfDWkFBqKURR3q32VM2YhbOh08R/v+Zk4tw0/cf9l4
uMqkDWq97DencMR6LyIsStF3tO62fDG2mFlMTnjSfaT3/rMXMegWkXmWBUNSqyjTeAxo0upWz84o
L5YZWfELKsBHcRE1vguZsQNCBhajbw8rVEKTU/rmSolJQm+PR1QBOOJpV5NEGXncyEWe/bydPAU7
Fc9gw952G1IIT6Qj1i+m+jzzJSA4K3RNnAFwpItqc9ZOEncQCeyrrtb8S7XrzY9XeH5EEeGA2eBU
Ozg1LoQbII6Z9Aapulzr91aLHN/zQQsVnBwhMo1B1AtneyfOwZlAt4s+13VxItahtQvnznZYTi5t
QuEQ016vVmTrkaS0AqvOuFpLwSYe1Uk+mqV27ZukXgBvyITTXb9eM1W0Kd49hLa0QsMYhKIiEBMJ
59tWGe32jm8QlO9KeBiPH7L67bpcWnUKin/Hp21MDBpHMnZEMNAaniNXZFCiEk1dYz3goe+E16UU
0SqhGVNCADR1JhzQUCevYuB017aNCuKlKcmuxcsNV84Nboe41nIFf2M0ZXpapdaKzsspO2ohPVx8
yV4nMQ2XKYQE1HNWeVHM/6eH2MpYBE4gsbYB8+sbjej5kxTpAYNADBOoT2yZc9A1dfvJYqCqmRma
ybac9wVhppSNwzksWlNvlVRwEvWfZDChuTZ/ryiqqWLGZyVCov6IACKwdGdVnUxlUJgc4VbX3dTo
/cbGqL12yKBvK/Fwa+Hst7ZMqQK+XJx3jOaLgqL8wZfsoLdEoOgqkIhXOMS0/u36OQOErlXTAA7L
PmiALgmjivq3aLPEPneUD0O3cAinPBArKdjkTbMxP43eMea1cmXXfJSsarunbJ4JGmfQpJZhdLCE
s6hMYF5iOtbN6aO+FJ60YkKwRRm64BpgTDLG2ZEXxD0+NbCf5Et/TDvjvIv6ds8E9nELhdVDc02p
TXEgTOp0p/xRXbpBVsUmKTrsgt4Om0CzLmyPjVFHIYWBWl4TFFC4u2jrm4gF2ooo4u9rxTtN7bH/
UkAuqIp5wbOXRIdZ4IYdChtltxLTyvpgNIxA9DPY71yDtqzwe8aRs534QJStycW06altIMlfMyoB
H2xqXUklfb7rimIQ3xI56LOI2H/kGNmAqQOd9SLTxL5OOBicaqaH2KN9UJ6gQSX/8Z5c3HBpbJGt
jIWCxXVuqK4r6Oqmg3P5u+nr/FLwDjsJI/TLklC1AMotrQKa0+GG2lBOGyev4++v2kku/oAtAMfs
trBSlnN82njHNYrT6tYRMQlEbdYPSPRa3e1hfc298Al9SN5IbqhoBQBNWHzZjPDJEBXOCCIuEur/
FfCN0RMN5V3M3WHd4FaZuVtcaJPG5pmbQrFvMoEs5UomUtbTvOdiTaqvrrkVeWFxjUolfGmI1NLA
yM/DoBcS8FaCNcOaYHS4k1DuKG7azES4KJYDEDsFUyAS0KYzNr0gU+EPg42GDzItqPrlYzEs1+6o
kzNmniEVXH2tjUjNQaNATlmwH1hk+H5LHEZzReLAhZMs5CnOpIuWZc9HEkX8mkf/nGSFYCXcDJFT
C/EfcyZMDfRQOI65K0QwrHlF9OMcvesGpZZDuGYPAU3lFd7M6v5ZTjo/coahFSzZx5f1hU4l7NAY
vH9Xr1l27+DMy8YLbVMm6NSRgI4SSKzlYcu/tq3JHovYuePszjrmHlGQjRU0GUokWcfAMO2WhNdq
S4drfHk8manimOQq2U5cpT4+WBk7ikDJaD+02BkfT5ahG+ZajKxXreQAiWDsSrCnI/QjZYYV9TTH
y0ig/+tfBFvNyzeaJqdcpX1vcuVIHUp0Gf16jRp9vrzKB5FchULencRbZqDhu2UhhIhLBjh8m7KM
L7gmvNxwmmRHPMLWrbbsY4/jK2HXczgFU+XSIKwhap03L/YkbWq9OUl38egj204MIdiZwwT240XN
GaZ5B4o7iXsOaGUhkYWJNt2US/b2Gt+ENIM8YfSMLFkPowPqQ9PYfBjrXeGoPAod1Er0nIWIMt/G
Og0U09C4sxL7ylmA9D1eDK6kCOYWf2KwvJsGb/5QiVaTHYTpV3cilynDKOdUMim0MNM6fb91pNSv
NY83JfROAkXTQ6HC+o9bSBRe2hqB9GUQ7BvLuvRZq19JUg0b/8nRuJqbOBsJ0FRS8s0/dF+0nEN+
VJit0481t9/O83DIbM4XehEB+YL8U6LYtHIiXun0MQsO1eIYNwItTO1u+0M14xfdwQBRPS7gaGpq
59arVG6heLSL07yPLj3heQodYLd5Zrh8BKKr6nvl+9HHQyxuMkaN/2E5EBBJM66TWm2Au74nxyor
G4ygT9KeowsofeBP9cPF2BOoTrox0aNYLqksI/rjcPPbj0UU5FQysrF4D04diquDeBDcvwlDaO9y
cBIq4RPtUJB5DD57uoXJwl2tRc8gws0ttrSWNYaJcoLfPh0DjfRWdbXw/kAxQxqSXHBeeKtY4++o
k/zwCdi/7f+yea5uhGO4UyfmLswxl/uv5AvwkFGLL5CqBYRaEnHqHHaO6TvY+LJbfj+HlT2copod
MnFSp7jaNwWG1QEsUYfJ566ZS/FBSt92t2au24V5GRMk0fPohISq4xEfBg/TOpCaikmzl2aj9LVh
ijURMp8ZUG9x5/S7Dl9ObklFJcTIn+Z4jc6sjwMTuF7L7K1dto70d4qX0/qja0JQfeoQEIjPELFE
pB+JaD6mTulfs1JDFPrmFCtX+UntZkpYLHZx30C/w50y2D46PIPhvxdovZZYnha73qJP84BT06NO
CgV4b3jL9PVh3Vdkd9gLmkWJIy4QHnMA7stwsoJp+InCm7rkUFHuMDmSqSRLPx9Nn5tjDLbYGKWT
2WS8koLvrxw3q3WSjsn5uagyPgYmZjcJ8ItU6X8r6C14WDfLW1+u/G4YUHdkXw8l720idC60qP8d
i8Abw1xPl4G0VT+zrcn9jKVkinCRWas4+T69sTihsjs6gdmqKPfmIvb7HJ3G2yWcKAvY5ltLUdW+
YYNi5gaxGM14RYV15DAOqbPnTP6Seo8SSVJ0RoPb7M33/B1m/knrsMPxhC3ejV+Kvf8vQRCtn0dY
5pYHix9XlwJzAge8Uqj7kLKIppWLAMvxQP2NSrrVCD4BW1pm3/Tsvgv0lxr9wlwQXy33zbm1lWmU
mfp3eDpi9I9iCwmI3bKmkIpZ0WLc19o1I3s1LjMOXKrMneN6oUsfADLWdq9R4AzJ2jTxurdYD8cE
Z5F9st+818JVow61eiGb9YGneMn85AYYMrD4i6Lj2scDuKrs/JsSIkZPe6cU6M5Hk1gA+wJtjpcv
5FX9kFB+uxjvCE7y+FZJxo1+sjmtl2C6mnu5k4tnJNWJ/d1HgaqBGdNyXVZ8bZZff7QOgv1H2R+A
5Vp1EcGLlDWTR5G75pDgkw5fbdcL/mvKUFxJFzchlaDV97aGRO9EgI05+HlFOi0yWtb1GTR46NbO
dXBysMKmKPtRxleF0tTfVgOHxl4fQ2z0MBaC4Lhj9E30igvUfMJ6xtHfQGy7WaEpXMyUgHQ7JLgk
wdXo7Zzpjo2C0jLSJvtKdLloGfa2u2NOSlpEYamwEEfo/1YITzT1g8QVTjDBinkyHUDxaMR+vFvP
1P3HynGYLn00Ys6UKC/uwwUg2R0ut9NTELtUYoZuFBwTqsccXv56lUgfmDUDdWcK6eHnJIrRVw2r
7vytJPf6ld0gbURpTSG/AZwFLG5XmRKLgaWiTtVub2D9KIZGrPmqnbfofpwrvyM0e+AqBMOTfr4S
wnHn742s+Ih5nImRFroCPyPqLF456eJz4QKntzi8XtYT5yqUsFzNeactAugn+A+N422pWHe8+LSS
k8nZLLkcF6I4nvrAf8JMmmo5jIftXqXMOetLNDfQbYP2bFXW8qRLZYJUaW/0HxgyzhpqN2fTIroc
gh6FjwMBKoLRXxXy9DbJL044Cdq1iyhFeY+s/mOo5kk5nq1d/df8DDQuF2SPBSgvSy8BySrU+aOr
epN8eRKORo9IlXu4B36pjW9CIKypvOVMLJ47yrGeFP3DJ85KVwmCO6SSqOMHxMAHpbzvkZUAf6Sx
36TChmjrB2Fx2ymNpxkJIS37EkjcP0Q8zF0U7qS5uszkn92umT0EaWEQRlwx0fUgUdXd8XNz3bFD
xLBX4yfOJ46ybr10zLXc7qZoaMEQYnpPxPgFaPaF86QLUQWmBLuCYBE9i2/Pq7a/jV0Nleu9ZgTf
pbJ+ARXyonOPpQpvwEHcs1b/d4KWtKgcjw2rwXQycEd7pXgY+U+pc7bsXBA8Nm+5OdWBYLpkGPWI
A14b0HF2uSnSn8V6RaQkuWLDqPba7fC5vV2YC8kLtROrYiq8Kiab0asbmzprlX6J1zn7sFod79gA
sCCXWaxhivy/XLUma9E/BAwbXYAu1bHB5hEWmdPWGJJ73kpkGEHqmZcRASh/0yolKgHZzHq+1S+G
iskEfVmQIzyqCTsEJGRkSLrZ1gHUPMSf/MPrNVRS7TmMbNz8ROOuDmIJ0gi9lxe8dracnhkHqDv+
T2lHH7Y2dEe6pnhVwj8nILrP23REHGRHi0incj7E5/jEYSRSyT2uk++AqPnvy81bXYeFBgu7eBON
OfSww80ngkoSnPnw2cnRfX88PTQpVUiqbZ2YGO+zoVNv7BLg/x6gOYT0UVI4BNP5sQS83kdTJxdd
qAUu/4X7y/5RM8U5/sGG73uORKIe+iWfH8PKBUtwl+heBbbJ5a1ZLFnKufoT8mirLA1ljwZBfp1U
44+5a7C23zMr7mCPg3oSBBDNfcQG1sKdK/OdBC3H15KrGxkKAI2q/8CishUZkLOUh52B4T1IpT5v
MytYw+5ottkbZMKgAF4pkvhfPuP1S2QSqNdvTHoQPyNkcgQVEbx6gvYmu+vtipcpsEK3kRwd74wH
Vb4Xl2+Mn1nbVWM5F5pSvHeCdUzG6hr/4sMcsCtQg3wtNkTZDfQ83/CYJ7G1i0xXIYyUy04HSLEy
7Vcp7LsoUJM380x+tEGgV5hKP0J0Yyrv3Of1eJU0tS/x82YLpIGOCbk4GAsmp7a8oX2WRrHr2fvl
/BUPwfsvrgXYsOrggSFaZqtsnxrFjLR4OIqCsZ3CYvHVudHghLNxQwhGwMgiBWfFlXxnFI8H2nAZ
BAGrek6Je9C2TTDlYSScjQzsIDSjJXdAxKbIyLRrt1+D/a20mI51O3IEPc7gDD6o1yPaQKRNf0c4
nFpzamtgUSqEw8AegFwQxxvbskj90kuKdmc7vT6tnu0O7pJ3644Ctxp7qQ1ItGDBi/M80jww6jEj
8TtJ1Uajc166BqzJ9jyimf7Cs7wZjZTfdDWsfkFWmuf270cFMdOIEp/AKvq+gvxIlM73GsaJs1Bf
+lZEyJyqJ8gaf3/wPoLuC6l4SThjLB6Yon/Nz0p5dhh/i7/8tiBwENw5pCFxGYVL8eJrqS3cKszA
pTZfzWUFG1veCxmHQtgJtMUlmYAWPNl4yt2eLL2TE7yUFZSzdVtrfyKbbq/6JWlqB2ZrOQBnajYW
MBTJbcI2exl//KZrZyqaW3vpN0BhpSXFohV4WGeMu/Aq0dm4qn7g59MO5VDK4Uy8e3anSip2Vwpy
Vy5PyavlryqkR15ckWxCyWPB9LU2BUGqbf519stM34vvi2PW+jRZ1sjWFWgkELxZSRqxbfSVYDMQ
iFwZV0Tf2OeU/F6dF1Lqd4MShLyAtAYWwfrwuIRAweUanloZCHLl+E1neRAc3umWZi+MnyJjXgKt
RyRXRmMjbfXKZRDfuNs926LWLKxxNdZcMaUMtwAD5LV6vnODGCqVVusfFaB1M0R0CKS7Qily5AMX
odhHlQRlWpdBe2Kl8c3VubO4LD4wRF2xpLRNZmGnTOtCLccNeo8EPAEwferu14AnptyDyLYvtRUN
lo2u1BHcUl7u0ovgrLkfhEZPCNy3uNXmkt/YwdVmMEiuyJ9AVamtDAKlJR2vNMhmVCFZwjzrihSJ
RGUNToRMPmRmeWSVpqVLvn4e/3ZNb3hN/SrHEaCLr8Rcxy8Opl2GsVMWPaLDz0uCQ0FDEq9OHEAm
BSdnhMg+09H7FRbfNAEZP2tAXv2rMAdP4lqQkh3AUWqZ2BzK1KVCsq/AOUV6Fb3A6movfdQ7YoE1
DU2N6t3p9k8Q/l9DKe4qrVyrJQ2gQGHJIWYIPj7goLT7OTDJbDf1lW6Cl2eqZsHk+Szee4IH2hqj
VCQyiO9i3ZA7MoQSVjO+XWb+Z3n3ZH0kMLzlqQESCjr4VHqScvQtBpeF4f016JYLA00jbEC/KJTF
BpOXo9qZOqLi4hfwj9W46YSpn/90GeyLhwojdNeXf3b7VNJvn9meUPIYT50vRPzoCf2jcyzDsoLu
6+rDet04HXTBy2p+EYZC8DpADFENd7lNZa6n7MdvtYhomD81QNPZaQ0atZpfLcfAucbiktC4qEKB
KKRo0eKb7yIUB4ZGE3JfpDBnb5ha6xVYSlo08WSpPQ13GZgM+exLr2VTo5XlLGGxn0kBJVg3sMcl
I8boP7iOr5UEG0ALipUF7u27FgKrs/c1AocEyZ1Gsu3jobqpI+THg+hnowzGt8u8kyFklmGkB1Ye
/+utnKDVKHGGIq5W9BQjaxyCvCX+yf3ZYztTRTnC/iHSjs8xXP2hSvUjmaJyNMYqh0V4zUHKGh5x
zl+6Dlxyez9E/Cc9gegxDbWFnzYuTrlmSWgp0j0A2WgG5tk6gOB2fggGZfFAU2ECbEmCCm8WkOIv
2gn9zydBZx549BNu6arwwEbkpxCN21IzZxWaFGDgnBBGwXmSfU7/UiNgW7XEUHlsfyYaDm9fR5NM
oNYS+PTBXDUR+GWbXZL26Pc17T20y8Iqi7Bctp1P9L+kztOmE5EM8l2TylWfrvi0jQ60ajotE8q+
YLZVrJ6beZZEivxLcuh6dujpfAh/nCejUieKcsYGkL22jiqEDXBwSQOHJbojbee1qcaguxIrnJiP
/ta0BKxLtE3pOzokLSFy/8hBlwZLT2apAVzNdylmwqQsVwVw+0xM8PPOO3AwKqt31FYvc29jWKds
HocOO8UL/CJzlpu0UXmI7mDDmS1dru7kfBzqD5nSEcFJq93cWPR5HbUoyXE9C1csl/wsHTQdksJK
TXOUgYlnF6kB+1ceTexvWiuCC6UNiLJcda8rCjLvClU0LRyRfRR9ljlSV50rMleK2t5jmzbK8z41
zYjvoG/KuLeDEr+i6VFm1hlI7muIAzijai3tViWc7T9D5nyzI/VIamtrmhsiqiSwmSdbadsp6/2F
NYOU07ToNBcDNHL2ErY86lZBneayQjrPI4oqgWVUp7GlII+6kF0RuLlg4ZODRNjLgG7pmMoqHPIu
CCdEGkOJ9kE7dxNLMFXBHH3p4ehRMJ3t0WFTnS+JsOASCkb2JOHohuFG0YzeD08aWzFECp4UdZ1J
wTJCXB2wWkzHegJ7QAWJp/27PxXXhC/PtcdbJVwszBdlng5xogz1Ij3qmDOgxuDKGl8ds4666RiM
WGjsZreSCKjs23smKBRdB9QInTOI3lrOQ6qGJNhbmZcYoS5fOyqazg4I8LudZteVAPZ1dClU8JwA
uo+VgSILluOj/3PC0EUwZuYIXKguQUReG3EzSv8v5p7rOxRrgLdcUdiQ8VbqsKBocRmD/LrMIlU0
xeh9rcjuu2CbtV+vst4hTLB7GdAEST5GnrGqhbj9FHx4i5IYda2qkQE6n/lSDT70F9HPYr77aWQU
BqKdO1g0bJ3Dvirh0NypPBFj8Ey6DWtWJssDW7mF2mlvaHlZVBmzpSN1+Dc4EqsgrTCR9kLbM+Xh
2gp4i0Z8o4ssFy6H3jQVjRuuPOh9rrOdA1BEuFxHiRizTwOLOsc1i4DbX1u0pR/h7ms3efSkbcZ+
zRFv+Dc3hRGYvuGsyVzkCXmVoAh0p92jYHRtMnBAUut6vbQATGEYGiFRvo5/erbnDF/dSZha9Acy
Zs/JR5YZ3g+R5S/8nbUknDwOqZhfsAVkzfcB/fi6D9J4EofUVpARKlJtSecWyWYblz81T/xeMiBT
z8RK72Sz7hMQk/MaE6jgLJb1wY24+tGuwQ5MNDNFZrGBAOocoH0MehL4eRAxhcPeZ2alhLOqqJ6E
JqOWBA6bbyxbadvXJ01B+e1FF+1z/HU3vqeqbU3LOkDj86okZiqzPzgZZ6njJY0LfG97FiqscaBt
PfHVEScbWHzHbtO5hU4H69VMw+wecisIVXc57YNQPjrdNvoJjooPVChF2xstxwm/axxoI+ZU03F0
2iJu1NIRH2R2EaR0sF5YvVuJfMS+Gi/gxlDytqgJINaPnT1NGPVlil3ds2bfi1nNJDDcn+62PzzP
5Xi/VH9G1VjNZpa4Yb+BprWkaoJ6WzFdz5sJupJxfjTutk8lArhkvT5cPPXP39wK/NNTU/2KexjX
4URBt5Toe18zQOKG0zOM63v70UwnhyqFvwK7JHh7iUT/6LC9vfHvuNIFhFfat6jEVB1D2iqniUqD
aj9tFyKEeBXvzLKLsroekW7WXs3nT94mK8pYNLVeplIvibODdMZkrs0qveobIOZOhdFu1sqR9GpX
NrL9BcpJGqZuIm5x5cX6EqoUfc+nbbc7AO50unG7F3dwIDrDZBTO18CF8VRueHoHgdQHRweMWje8
KcxQ6Au3gUTD9ren9SGKxgmDAhFKIPSQs2MZpU5W3oB/t7obLJdHqEno4uSBpvSl6CUZEEVAatzT
sZl2/M6hjO0WBPIicsq6ObLp34L3FgF3Er9NJ5cEY/DfRROCOIquVj6BwkHsBM4PuJnZsmI426FW
VaqMCGQB9RldzBctEG14fXVd/wjcUCxbOWMCMvNu3aBkvXw5dYv4aYVVnN+7sNfUPYmZPJ17bLKs
qmBDiIJXAT6lfbGgyJfmKcVFosR72KiXPpdnbrJKvTaI1/fTpoi082msqfiJ5XxtlTdqX7PYMRnq
09V+bzgc4WV3nSikdi1AVxx+fFeMSX3UyyT87zzcNTpGYJWrlMulfBvw0QpEAC/mr2viBdogO49C
SW+TRwi3FHVELXQN/R0O9QLvwQVL7EHCYgqRnwwXPMWSBKWqbgZo4avwESEABGhGwvSHfE+Pe/rl
vk8uLSfGX8JhBFo0Me66qEUrilgdrshV4ogphV+lskKED8cq/sLuVCYMaKVk1U4wRlCWbnxnb6us
UHbMzvAbvyF2g/J24WixY4MJOOvp4zphx+quic8/76CbciP3daqksbj0Edd8LBhpGmW+POeOcnSG
IjGpe10e6aOkTTDj2TGIFmwJvJqT0PwQphdZndzicm9TTajOiAHqu4/Gq5URNM8oRAO9a1bbsNYy
MgtCxe47N2CIkKqQjjIArl+frlLPDRRVecfI8xeMv0jiWCdalwUnReRXFsrCUEMpmBVoCIrzfC3F
Rn4YvWFqWny++c3YLqbY94Nm69uO8pUD+unWgdfcOI3ulpaXXCRpUZ2rpZvo4kD1c8uP7B/Zp1zg
+2KkNcI9gIyti5C5f0P82czZDtK/ItkG3SxYhJaSyGY/REjoqKZNbDFYXm6Fo6J1fAE1uHH8fKlE
Yaznq4867T1GDib9pj5neUx4fpweZpgG2H4iO/KIUvm+SmKIx5JCgSiUIZOQyFtW8zss8QIurDK9
j0LUlrGzX4O8ugsNJSWn7FogZ+esAfoe2gMYwWdAkXPbUdl4y3LLGYLsOBEbWYy4QSFhEHYtzWwv
WXdyST0Rqgy/rv1rwA2nP7clY4gcoRbcYWyvkOEEccAyPk6zqMyRNr9lR5rvWAgIlYiRpEshl/Mk
OK9K+PdFV+fWTWjNQXbg2A8XnF5fAsCeyj+VaPiHkQx/pzmwZtla+CHeRTjDFrF4iuZxkFhKYZ58
Xwh2AzY0eWshY7Bt1CPBRCKX/h+rwM09Yzc6tEpOwIP32zRlXoYp9bAq71kCIHQCsrL98JPZ38Wn
NLkzWrM4JFJnfGHLTAUDgYArb1+JQ5OJ60IR4pRfb0qErOaGedY4PWvvtfKUOyXGRoRwW/xRQ9EJ
Qt0aHmjJRkUD41BVlh1zZAz4VxXHSnc/acSCmx4nPOhid3CUxdS9f2ZJ6pkDsHHq+1pn26CiUVhm
i0olNo0bsFROxtj0hyhQ9OL0L7TT73UG1NIiNHE1rxNmZR/CNK4GNW2n6nR1Dd+kRkqnNtHZ3yc+
/2L4dthkKhOr+c0E9AnllqDxwu16ppRdXnVma03CL8JNGT8urfHe2NoW0Rf/apfI9ChphghdhyyL
UTeGsqGDazcxCJdgsfRbjp73+MLuESXL6lhleUKmmDyU4VJJ6eJi8PgLn8JeITna6oNFvdDImzOi
gMBXTkhXAm0ygSuo7DxTwnNmK2waFYe9oohWWEX7IlYSaVwzEWQdQCjJeSt94x0jWGxJp1NxbZte
Orpu21uspDP2TQbFU7hJxbuNzmyTcXyboEMpUqOwXl5izWYmi11jh4cwLZ4t8VFRk4KMwR/2xnu6
74BXFN0RcHYw8bkZ141nBU6e7EgPKSISJkcqzzRotAetXDntlF1ejH0w/lBppzmWmzJtGnrSqCYx
wuD9ZWy8tpjx7lRDxgd6zIyNDEu45ibnTf08iIQrABksSVb5q9nlWQ24d9uVTiSMKMVyyuv9ihS9
NwTa7JrEBNKmgCym201xb6+f2CnYSOSb2ilSh98F5H+ztku9fQpqN+nbLh0kuwQFVaiSoGoOeSzU
jiYTmQf1voQm84+nVi1Hbz3htJP0hLQXJ+HsxQtlZKth+G0NfDQppBx7JpVF3mYRXB7uhVugHIxN
+3tZZ1+5WpgMmd9rTfCMx5nJtHzQIutcVGntqvUkehOC/GwCpFS2+Dn++M9m/kNvuqtuR9ur9N/g
LbdvwfWAq5MJHBFHjVQscRymkqbgTICVIp8UJnr5WCgiRqhm52wdI3iGS2ezRr1SdgK3DP8aQ091
4DMzB+F9QZhhgZAnKHI1Nrgf+Zbbv9y/W2ZBKywcprPNSMJFXNAbfDxJ3rCiJoQ/nyOPmean5Qhs
K7uV0kYBNTR7a56MXQEW1voCtZu1hTFgKIY1cOpeUCALFthclrDJABmbyJWgV6SrbD22XyGGs/j/
T54kSKImOjkzcC0toybcgBaemMvH+IwIUer9U1z51eNf9PJzXnhRWuQgpeAGE5oEJeB9PLYCuLJM
LaUHu9wKkSYRVLZ2ncQKV0uH4cGetDQinOaxqPrz6ZFNUaoMoY/k3t5xZBVrSkI9lCWf8eG8fon9
Z1pvI0YPZlID4yZX2+Qdourkr0BVbfgnSTC+U1EVBer1pPuxRnPE0D4ju2eema6he2e3XJwEYPvt
Hk8sLBC464vOkbGnUtt3/QjMgyZbClLMBWopfNGXNkDqS45AGAbFZK9eYNCWQ8LdScpXY7PFueIu
QXh1cNgxrmOaQe5iHykvo4/FHInH7muttPIZxBkLi3NJlhzaMorepkpWTqloUhTny4yKBnHYtp/U
mXZIfWB2Zij26+UNIZNQYy7wiSHmJGmjEXU2YM+CQtg/vjgBniU3EviBAMSfHeUfJTHI1O+4TWpY
80zuRsWoYIaqsntIjsJKvhnqD9fTczPDFPVRJC47pXQNdxiFd59AbuGuxjCUX6/hzncB/beodb+d
feuZBsRZRyMQ1mO0ZPklvHLtCTVxjxY2IcUEzJe/FrD9mu/1cgzZhhX4atWYfXC/KJmLd1MFWZ2y
daCh7M0TRjyUpEr6mXy1CYffT957yIXJNFYPZinD99YAbXCb1786hRf19Shea8VMuYccFupiwmDZ
+2q21Tt/3pSml2/5zHpQC+tu0VYu7tbs2RaXb8wT6GFqnvlHA/2HLIauLuzs/NkcKaLfx8sfJZQw
TF6v04Nn/OHTNV8Cf4HbxcwnyS06apc/zr1koxA0DjVruyMRd6+IfpN2Wjr0qHRkBz+g0V2gACwc
MR5ubG6SpHO2RzTHJrMxid/bViDod5BRzBBNf+hPSXeGFj8//wIsSWEWG9ga8LifCcHwHeEIkihK
8vUG0o/H3tyvfFEPja5gNu5h9N5LbR9JWMkz/O+N8tY6JdguFt8dsMM4DHHKJ85AzWeSetBJoTN2
FSQYtkiW6ei3pgcw7seD1pcVwOoa/EK/lQtH590LNXRmW2WDbw+ncru2+frtMWDlOK58Wz4v4usu
sbgOOzCYCIsDgyQJ6HLS6fYWuOauPkiKjCx6qDuPp3oh3hka5HsFDO9/St2LuxD5ABBanBiouq6r
jRyJ9IGf6bw+wLogyfYb/KnB5+hsKM5jJcd0y63TfSDYTwSHC0SXrfthElfuoCgBDR0ej08XljkM
TDt518FoHfZlX1tQASXf7bIkjzlUlQcBpREO3SYDV/iZWuUXp5jDhAfzcvAmqiJp6jDkmMCmeMR7
N2zsxAem3gFb1S5wy67AdTuYoqsp/dqq68J3uh9OjzDyLZyOm7JpPTniFGk64tLp2RUHA97m4MD/
VYs0wxZMlKgO6i2Hvpucg4HJDzFWd9iXPgQLEY06c9XnfItju/A9LG1gmW992VnJAMq33U7V0+hr
clt57yTCKZTaYKhKoxqfDSOt9yhoIP/jefKH/WPflWTwCrJnqERofdUoUR5ExiB4/B6yKl38VSdJ
sVJUDexaRjgBI8uAX84WxUHdWvFtnjHkvdcuoUJImz299JsaxOSFOEWzOY3c9NBsioGylmjp3TFQ
N9TgLuEvCefgDZd+E2qJimYoKjsZvtATafn3L6s69lnGehoLDZApE4DVlS9Vn1t8GN3mtRuhU7E7
qAaAs0CFxzM1M9Mt2tkRbbCYxJPggkmwFKRMGspBHECi3wLfQWOcGSXdmDEXr7Zg0KJdzkLsLAH0
f6LlbDBAlgAjdOIRk9gCvvH7II3ldNEMYk1e2Ef7h6df67gUbjbbWI/9z7aAofPTKSAKg3HaBGMp
yyYePYijXaCPOQOMHNJWUAzHHD7KeQqxamOsaFzOEuYt7DE8EhrrgrJD0UDX7M0ML4yV2QQf3b+i
BjNahvgnqM6pyuK+GhXT/deX9FwwOfmqTUI7C3KNPOtEf/ELU3hbHvW2XM2vkIjt2ms3ubgGTZFQ
OSbPZ1cTTYVVhWvigJ+jl90ZyAWzU/T700QHZuQnTF2g2QYp7bPN53c/UAg7HEb3QEhh1C9Iwj2Y
NQRJqpIOWNCui1rILM8DzSV9OjCzpYa/b1/9SaS+ewrN5cbiMYOebZalEU85NWBQOh3Prm59GC7C
5jMPGhsK5rEyP9z1VCjm6Y3Z28w/Y8B+u+Az5fi3k0rNfr60vsTCO2t0JC6twxxvRM8xeXtQrSCd
2r+U9/uhUvohVYUBaxuhYeeJT8QPswCmJI2YhQMSzTfHW3nL6oHpqsDOYFCnnFWE+IkAIxlPn7rC
Iq+Qdb8lF9YlORrHmG00XDPE1gBdsA0QCvIDQmYlZybR0TgYR6FNowJChpqnISuUXsCFZJABPR9W
b/8QEUWfd2wd3E0PeDtysj39WggPd+tbORhaWZu83dCHBP2FNZ3eewFbRwA3o8U8uGSPsI9X0rK2
GpDBXUKTD6pXUbzMlQrmrtQ4Y/vqErXA+sOrxJmHS6gAvkEXih6wvbuKZZGDGJ9Df+pmCrJUD9ry
6cJibsnKXdAsZSFpg/eNWFXuy58BkX8jctWUrple9Y/34nifIBdsuU0Ye0RstYSwo7u2hxndgnIa
jPPfkBxwIbhj1xdVnMPf4qD07WrHc1MtYZCG9TJmqSHd9kB4JMBrDgbU2+ij+u2vS5DeMGqrX/pa
UfPoG9rzQo3z8Fabh2XfxEFNHckiPCBvjpaqYUiEyFUkKGu4zqY28WgHKa5k/CTV+FTRVPT2tBTd
6Oc+/UWtviH+jNq5sc/lKj528ttm0vKTK3yZiAMLhaV4C0RfG7Fc5S8YAQh0Th7X6nUY+PDAwreG
2JIIu+3PO3gAeMlcD1LBlJ23nr2T0uRzLt2O34VTpZ77V5pYbrUHB/am924PsQz5F/bJWpL92kL+
rBZdD6R9/clc4fJAb6d0q2fT4eXx83xrwk5dNDNTbVMuWhkOcb2hXE6Lb6WsP4evMDOmdWZzUdCC
79P3cTJpE+HqqJK7GswXUk0gcCwpllR/p57MrnjXVJN/DtRqXY4riTvdQlPHRv2x2YEG6kKxqwyA
d3nh5VOsKW87rdREwvKSaRrn9q6HRZyA4L24hzco0hldfnaiqlUOtJWjGBi8iHV6cpFt7DMsF9sH
Tbhxf8SxHS1Vsw2Ch37l8UzNHlYlaH0Mttl6yVNe0Gugug8CsivoyXZXw0U/y+OnNHQL/hiCEPES
HU4/0e4MTtf60PpX0hPD0AzwJakFCD2EG7KiD4YtzlULx6k2g6yoXRrxs7PxeSc0dptu/QGhHmcC
K6XtMs0leNCE9gR9++YiOHMBy3QqbX7AcP6cqjZ7RncGrh+fsijz/FJ985FBp6DhAoVrSs14JUes
p21sl8PHpdhIpDuq/jCNA3MZDif+f7OCnztyr86WuehjWAYBCPKss5RLau/s/4PBruIme26kTt4K
TXFPG/tQDPgzTV7gqEzz5UoZKycq8+8lcWY1UjCmGOKMEGRXA1ZuNWqYgK25qYfPiVDfhG44P0jI
NPdF0XJRdEE+JZFEaztOK5MPRXA95VCvl/rxpUOLLncalKCFw0SYCJs0NPC+e+UhwF6V85Wipchd
cAx8h4/lPBzH/wY/Bx12rA5WFprZ2cz65WBQBgbRRVdADVYOPg7/glcNHXC9iQv3zUWcnP7cXABM
CUzYdqMwA3A3LbbjQ6yG28uz04Qk5bQ4JnP2vYze07HJ35F0A2FsRQVNlzjzMKIfxrIYTDHTlNOC
OcZDEjNiJxR1lhI2iW+FEEFZApUF8GIA93ZUCSWP2aXXqtVPXoyxikqST72a81TXlX14x7qEGt2I
n9r9QQu+GVkGI7+EEjWUXlZpTWEzKQlArfAC6oqvHYPnFrjuZZdWstOpxyS5KmyZFxVIZAk01+IH
dfSeqfF2xDtJH1H9bYyW9wOqfzEqORE/7rtCj1y5EemmLfWWRkIuaADeFLzVNfXPOBWXRw4yxtkT
5YzbAGSGobXSkqsrzJfxAxcm48iRdTpMMe0d1DY9MJKMazjxU515ffaq4THVzZNizbRtttvK84Rp
m9g7h2tEkzzZ88WjMgV3nhjjZQLgVIhwPmEZqRSZUroVF5g++4Z+bpaMPEkrZwtpEI4QXwB7IuDX
RZAHVBvQCQYulKo/EQND1CaIQLqjZwMhSyhKaQPFtmfzi2cpiP87u2M40qFQ+l0KXIhTMuJOWYhI
2AYi+wg2cY8C8TKKCBLRrqsf1ugFWsFPP5Ir7CFeLdMjsxSAbYQHLfkbboDS2gJrVA/sfAXiX2u4
bkSQNuqpnmZ3T6FHn44cwNWGXgwrrlH/dvDOnrf5jB1KzMsYznuerng5i92ipn4FKbZ44YKkx6SZ
sYgmA7NIiiwl8nsG8L0gcOtcKRj0/ix6O21AHkaTFpLZiliLlKf/8HxIWaVLZUAHDv2Oh6ltVfhO
yt7lYmrkxy815/k3SjrkaCgOyQlIeVoWihzKZJxaMjbassLf17y3U7n7hruvzhy9/QWIwrremBgB
0qruufeymgu/ICnpJx7cODSHdZjbf7Z5PfiZbJqgd8uRsX7sGvH81iez4+5qG213IgFS8Vq4+4VN
tp/f87z8suxNzuy/ZX5adVzs/MPu9tlEKaKvs8BWMWuHbLQDg27ZUbLe7aNm0RDtSperzHlKd5Im
wzyMiwtF7BavZ4kEevSMSjsSoLEHkddPN0V25XxRUwOtocBJ7GWrHS1zN8rlzoOx53vIgXIw0rDa
GXL0HM4NSSqmBvWmvGTH9jj7m6J0RKQnGUhiP8P/P5BuxhIlBr3FyFIzsGpIWpRXnVfNGxHKV9Dt
7/a3qCOOZ6q+kUq6QQBZ8vJ4z203VSplGxZlaXU9M08LXQjbpIY5RpRvf841mLv1ik+SX0o69/32
hDxYaPxcVNmsNdJkOsXEalUTCJZIk1TyYolBFuYaV4wb9zpWSno5G7qZwrxkrUajoefuTC5+cSji
ZfS4vDxZXDtQ0eJUGGQCfTmfASzt5sLAaiNK4BgWX+hJU2oULrJTVql2fM+ADwJ9JUD+H+IQ6A33
9cil5uAryUuq6N/HFLKZkcCB77Hil/LUxLkvGkaLXIM6qfGOFQzoy8Q+kOrJi8NzlHkQMqNTlKRj
kEL6ghGIjcTH36s5e9YDvN7FHU6vprVDtnLj9fqBUm0q9JvGGDMaPrrA1GRdnJrxyEbvqTds9Azr
UV0CrcKpfuiX4OuoR3L9lb5ZUKqy5MYYTn08AxlIGMyJApG7U1iHgKhGfx8zSOYOUMcPFN6ROrw6
U/Bx/1bfkqYyU8LV2iK/JCFtPhZzbs+eduMrnhTpXPevfB8Km2pk6T77b1IQOrS+HxLWMN17mVbT
ITSrTiTlL4eo67wIZmI0cgnwwmFwMoDMRJOWUxuODGo5r8X9bnVq1NiTT8SkxPhJSWLjFI7RWXiF
pUMzxBcDFMxUOoLY9tyz5t4RA+Tq5ifrj+MnPppIDwd24Nes2955EktoPATVZ4NL1zNAgLKQ9b56
rTLZ5pfY0AbB1SPn2kklg9uUxPXYZFd0kvXj3GzZoHIHY0pQQ6h+mk+OdeqWlAIfW+HD4Kg627Up
csWf6FeSYh88/qdPxa06z/TIjwB99lpeoVXbXfy8Aqr9FrJ09xFMTCKsIvT7lamNM30OapOvL7eI
75rks7VnKMJcwM8Sx3MaNx9J1YWgJ0in4BHAo5Q5LHDkT98/TiJElRz3xHtM21t3tGJ4Xv9jyzhs
kh01WQIzwL7lqu/jMmHTJBXkrJhUrQW+E20jAXCXDdeZN4wET8P7lOHlCfKDkzR8bx8wh0+WPwOf
BNEUR4ckLT7q1MnbLSrbfzxDi3ec4O17UPOkjPOUf3U6mL7SVWwEyKBLytgaWlh8dgUoOVtryebb
GdMFCv9k2+rHPnamHAuYqHSSqDjYLHXVJVxocwGQN6NQ+QWVH4Rt8xf/9Zp1abXyHZgMb8qlty7y
QE5kCwUR1BO+eNwq2IBBJggGdxoQNllbxZ8b3yzdaLL0XyEJqZI3Yy8t3Pw1S1yJher9L/G/rmIi
XrYDGsigf4oifVXC5BSFlnZeWbHqZM2S7NoUQ+7MUJDnnvCmGSm/XEoovVbJ3kgzZUDHY8E4PpHy
ixgIr6YpEPVbZj03yJdYL1FXVcupsydShFNKAie8ZIPlZEkgsRIgffYZ4IKUt6PwUP3+GoBUq3PP
jU/n+4h4KXvOdP1RMzVVcN9V+h5hF1NF0OtIXaA5AT0x2sA71UIf6nFsFDKANO+DeJflfaD9+RIU
Ml+Ee0QBFnbRJ73P8AtBKUyHTBZSUn0Dna7dxPUgN7uFbNBXFcaCqDzGRuvZB0xFdj4W7MRD/XY0
B7PIZ8j2akCWiIOBw3/gDUWpWMAl3MU5A/KiypiI7srfO57S+XnWuWO+fPu8XW/BCdWs7pJ5GjnZ
GInNgS9mL+ZhhFXP4EtHFxeu7wmBB9CEvfCexbi/DHL20oK5OYAtwiH5QgoxOh3TjF/vfiM2sStP
ADjj2WVq/oZyt+c8QAXx2XcyZgcHKYwZdHx7r7+BBiQ6uTPUfl0hB1KV6VrKIyfxVktIcIa2uHfk
Nj3jEz/m5tprCs51R9qDOEV88TTX/TLlH529RmHDYFg0gRM26FymEtg2O2qkmvgQucniCrsk/uYF
r8hjhuOqfrui5ZcKcw6VuWwmF1JrIMrdYI52PuwidQs8Yloq0LF1gzwJfhH+sQi/xIkEj/RQPzxD
V1NeSaeu0/FQ0Q2lb05bXEqoz+D7e4roZHAHCygdRxmuhD1aIJ8M5+51zUP+Cy68frwoDF9KXoYl
L5PFCKRy4yXU0bSJT2Kd6AxvB0FFyb1MWvHOFgPAbX8S2TrwxosWoyczrgtnnX0AenD8gcsE/XTU
ba6TYlNUl7zSiUVR1qGaBBsjJRYsk2zQ2SnWqX61meL3dLat7gD5rW61Ofvrs/5tEkP6yul1oVyl
b8701wFF2KfX194nmWcHYThzLGS9tVvkAVi9FDyroB7OkNJq1FuxLYIdz/g0w7pBj5UOXAIe3Df0
/hAXvB8q2AHZuJiq/oYiuv5AXxAE207pNyaa30K4w34E/1Euh8l+CRTyf75cDwHVjjJ+P9IfOSeH
gxOivfoNNSMynfh95Iap+BBwTn8b+BemxbzAxsVXV1mx31ILWx0HihfyF0+J/+/hNYgbubzKx15N
IYoexIl7dKSsFDeKXZgO0ZrKJZim+1OUWuTa5y9Xh1MWabwK8B7c1vDjFtMNPithGdwkEvBOoWva
+2VkDTdaQ4eAPmHUnJsO45OPvIkPgKl9sd3wAaRCNhBRXbf9f1IA6QPkCdS0pk/PvHDVprksDH4d
ABeGcts59eMYVwdG5WuESKPJ070HreKWRCMdHXIVrbzikYJTEh8x2KmrWG5PQcLXAtsFXRzPmv+3
bLHkumNeB4ZTSWGgFesYCmllq5Pna0O7P85T0HVnpPPdt+Mobi34kRjevgMiRo8I4OeC5QI0nNa9
Wr61vqMC1G0I/wwJpRnsdC5p7M7TpAUtQeCGzwHei3Phnnq4pVkY5LjwfTrweO3galcccI1azq+c
qVjEYHEoyY6i5I4w/YQMGU4ipGC8sZAM/i3Iriay3MMcZV7hSY7r4JSxvEbYRPpmc3ip33H4YrZo
p770SpU0c8EGvGRiMaRgRvh5jGCL+3E1XB1KPwgm+dXYfgGt9m8T+hPuwPc+bikrD8whtryxWu4e
IU8W6NUheuyS4Fkf1g1aHBxBBaeH+SFc6RPPJFON+7udMquUDbto7xlyIR1jYonL9ON8ZMdvGsaL
zeOqgGyf2prBeiuQA3ekT88mThtcD7O9z4PBK3J+7fXMvjpwBnm6pQg8jek5qWEXF0rhHeN7Vllw
+mxUazTNs8gnIOQfz0TVUtkehVJMPWG/eKdu+7dNo35z+HUJ67Pk4aBTSHNJVM3RLvZZnubG7C9B
DfHKrw2EIdjZn79cDL4wNoUtvAFlF3AFBSRZj7KVvv9xK5HaWSziPkjPXm6hNTSqi39hdQaRv076
BJ0ezoL78ICu5NGu/wutlBtmhvA5ijdcxZbRrvkGD0Vlpg6BI4GVBpq0ZWpYhv3zleaUixde+MvC
y1TbuuF+qD3FNlM4rj0Pg2VqycoSUahzqpqU86xmvafcaqbjcLB/RBS3FLHdfZ/Gjvl8F/lZepsv
opb2sm8k49v4Qate9uUYKJYo3zXYmM1a7rZPHHqIYHaeLWSzQZRbYye5SylMzSQJxkGtgKvijg1C
VbEFLiujU+g5bBtWmFl3/5PRgqmeI7w/4WrvlxBaGWHeFPePpAA/WGQ//HR1sBdgOOvO0KY7Qrao
AX06TGy5K3zV4wyhXyFp3AlO1dGhqiFcys35ErxfTz/6lcYY7iGnNqWTjqJ/gUrIQ6d+euD1QY/n
1WnmPegapsdSqb7gkJ/3PPRhlX0Z6+hrceI1vvpmwMErEpkq8ux05ZU1F1ag30fHBgP9wdJPpZDv
Hlc2+FLrDAb/EEwHxTvq2XlNBSXAZKD0q7lMphCtVXesxGoAlFeocWIZdNG1AaxZWM844M2XEMSj
BXCeZv0Ag4e4HeRYrhi6N1q7ZaIScTA0C90Mj60zTKexKLF7FEhzjFRFVNgCxxU9niYmc0Iq4Dno
uU2SEW2D8BdPPUZiRfofGaTydGodGwQd919qpVwv43H2IWZnLBVnEpjS9/yBmoGEeze44rU22x1b
TMATKqvGCCACqsjMVuNn8XTFdJTMAqdX5H92x3nEmPFGCMGqglEWkjOeAYLdo3IAZ+Oxpu6kgnVb
6fiDQdL7lN519com00Z5Z6JgooyvBjxIVaa1VG3qwfI676GgZO2xIF+n14Vaaqcu9ygAcXFGYm0P
E6MI4MRh/frsPcyX4mPnWCfNDyfDEkVHe0v0eLU3HcecyI8oubXRpXT2Zc/L2yjw9Wysz7m/nJjL
Q56RD+oyGcptmkmRfaOmNkNOgU5lxN3TeN6t+NWue1dTIMK4syXVUwtL0dOmJmsaqSEMvLM1ekqB
G9ZbNVTYSVSk8iOE//6TDxnU25yr8cLkZHmNEuY/DlTemyX+XO1VFUUWBoQCB58vBltOA0GffR5U
qXhPwfPbJvSTJb/V9XBrhyWA4QAgGgxLOKV3/UDEJ3WLg5wg5AxEw577Ck/nNK2vrbhEkUXYWuq0
kih0dW9sxI+z5Ou3OdP7VQ38qNkW529Rywc5ymdDsQhDHALwYX3SnNKM4EpNFTwlkkpd03p+4A4x
hpPZAM+5d9Kvv+xI7hq1hkmjp63e3iAf5JSH3Hv54va5DQZCFOnWUuEd6QQYz3R0JRfpWpv8oaA4
sywNyDV+HGoVgppwe6QgtDF3VVmxDslf457Qy8npaEzfKL5ibOr5jVlNqirxFkjWVrehaCmVIT9u
CDRpDi67y4jd11MH/SW7BJKpYkWAIvWZdeSadc03aD119RleYDGxfTMMYixxZK6IPUk08LeaiJUG
a7VkdM7E0FHM8dvFMxPY3uATSkQXGElu/pgcyye+yUBa1U1SJ3n1gcQMvpESJoD+x1wwRJIG8z3P
l/aW/bYNXsBIeboRvEujAYA4EQ3O8R1rJ0LI9WZD/OicbjRzNJch5iU2sqmKzIksPcxo12jUErYC
x5BdCPqZFSswKMkku6bdG8FrF86Xr9hi59I+4AkFWdToNbECSElA9jkVHAipU4Y0WAfkOGl8BpnM
6BbUGwfdlM+SAuq8d9Euzknr5eoJJanlusnUK6QQjxHmbZC2oJl2rd3gY2ozX/AbMsMAdq802dFC
3OqPrkWMiLmwx6hHB64KUKsRDqZWA3E76gU2WFMj46mLP5tEH6e/XKAB1sqryL5oojFL6M7Gpbpl
1Zp0QdOKXzG8+bJ5pYGrsyX9LVXKPb0or4q1MMM/suavM1z6rBLi6BDDyoQbVOPaiS7C2u0glcfm
eB6WReNZzbtoOVIvrn4CfpItqCvfe6aX4GGu5Q2Qtdcoo42fryLWswSuEv9x0KLx2FTORMqTf7Jm
VU1QxrxyicmvZZtw/vI1RBtKpibT1CaaSzmGRNVZ4syqlCR+40LC3tWln5BGpPIhkINPZ7ri2onF
99EsgL4KgkoVQAgtnqCzxyewHdr/42XX+K/0e+g//bK79xTdb0RsXPjLiiZ7yAArui9/4NACx9Yy
9cs/sB7wTZDRCaNmL2itKFRjx7HZnM4Cg38Kzw+WnVvMFeMU25Yi61cdpQ8WnrGiCzcM3RMBMSMd
e40zzPoPI2OEGZ7V+5JlvCwG+TYoSBqO/PutAlPtg247JGF8VeeUTwTqY/p1+CWGFGFGLOo5D/9+
3y22WEgFghM02vPJaRfMnVz5YNswLSrWhMQzTlK/nLce4rUCMI+/4+5zSDw1fxDWgeEeMeqLoJlK
MGNgHRIK/EJv21+xsbRlPomdr8ZtzeziNQv7QPcvKDL9pfE4CpSP7DgiAmlaiVEBKrTlwzD3DgQg
vcduZ/0bELDM7detsQZnroPhmVorFPkZ35zKUJasi5UcbzWDmhpZEroMqLAXc/fqs2A9fLFriV+I
nNz9P7/6Tpn7UN49EEO2zZpl4z80Hzg+jSovsIpdDyPHPU83KoU3B/Wm3nCAm0p7E6UYdwUU/tBe
T1F+q1nweSdR4px6BDwsZ/ThHxtVuiBjEKLE3I4eVAdo3NJaaNQbXQA6fcRvmxspy6LnfIUmzxu7
wioiRdwZPTukZb7UsQShpQC7fJMzmn9zcj2QWi0u/oC6Y0foAv3+G/7JSe+PrQlUvroC+4+/t0it
t1XbYPDi8ic1IGUjnY2iuMI+Uu6Pv9ParDkA4AfVPSnW2TlJjbMnOMbLu0d68tJpK83JIscfiC61
GSd6Z1t++mDOaehZc0pnOAp/wyJKW5D4sRhR0MmokH1rStAA27GRxD7Pq98ejiOO4T7h8DgjS96K
YRUxqkxRlDHvwclUkElB79Jhix6z9gi9B/Vqoag3n8n6Qcnq1xd2lsXor/kYHul+oVb0zoCiKjY7
yjGVvE1LhljFrAmUgK9TEffLOYSoY0LFSIrei+5d0OM5r+Gf2Bav++UOdVsfzLy6y/u0mk1hq45c
Uz5eBBYJFAxIkg1TtfO4dEoarmNDxgQmgmUdcbM+cD85HgYFjpXRoYfkS4BOPylhmH15htpqcCCY
URD6M8iZgjmslsGcuoDBGKt73p7MZosACQtBZYqiMu54g85djMiWT138orzk2U57oQ+cqSKijZTC
hFMOOKWhqlI040QlHuSMHGlvbQMJbdcw8n2i/XJZkQeFOUnNn0vnF/gFJ+y15k9JxcYCF12JqaA3
QNZSXtc2QBD4AyuSW1wWk5IQ/bCoFAx7eO34wI+LNY0JBGxONQmznSI3m02hpkN3mb5JmmYoLdl4
4V7zt3cHw8Zpy/GwL9VdXEYrh1+BCV/Jfxqw6iYTOsMZVMbouzvzDg+q7ofDRlkQ6FE2PsTC7n+d
GV2ePcwPphBY8WeT1QTTPsHo1IyZUtQin6KpjzFWiRGUYsXF/33iRzgo4UHYuynAsNDWAFjLaJGU
8kRYEN3LTBuUhwcAVqZ/DAG6CYlm5j/NACWIsB3vIhuTC4xSZL9RsSfMSvYMzZ0E3HDZBDndobll
3pWafacwrynJX9M/uC8PusAN27hutsSeTkZtL0vY0l4WeV0r6YjiVqld6mDJKwQ88y61v5Zmsk3D
d8o3RC2CkDothgzlsmsfHkCMGgVumQsjKNB6ExsYV5Q5xaNWrzJ9dLfp6ZtpNAu6SHAcqsEb3DDf
nDtr4YIJpk4yXVVjWo3f+fmnsq/dLNUwhjNiZGCarMHO8dqdWNUgPS2QiGeYeSkrnql3KPh47L8s
LOpXDNG5x9dsGlAFBW4cF40k6vT36faDAA30w2vhLnp6xU/DaBTRP73TLKXX7kjyekRgpvjIWo7c
6QoDNmaY5YUyQwQmy3jBUWD/JRogKNeiI32X1rmR82KlvFh8whn2hPdjgEL44fhCxrH1y6dCudRt
bdXm4tz0PVc2b22e7c0xpSizKMouSNn+Go3DimVAiBTMgtnTQvH4MaW+a6pkizURFV6cRheoaB0k
dY68A8x7tmSQzODI7YuaayUod00xvthDzJ1Yk+/q/L4Rs41xvnhbSWYpGmZ5DRKZRblQoqTqJV4P
6FAkrdfbXfTxuvHHzsZP9eTEQo5LgbUayvtheeXVN3fT+xYbO7tETeNk4uykqswpDnkxRPOAeWtr
ZDSKNBd2o/9mEuvuY23AA9skDjr7NecKCONO6sCxQVh8HCCRGmTwGDMRYBwCAopIhEXisSBKeFhV
ZoCUyVqItg6POlmC9BGUtT4bO2MItfL0+/uORet9YdOfwX0f8WjLymH9B7yGHsBGoO25psHeoem7
n+JbEwMqjM8lOeiYvEObSbp/+zZQUHgkh8AePpNj5dv+5pl/4Nzws6D/I4xPFNNSDzS1zHcrM3Ep
AU6FtL9PA6nk2UM0h4kO7EohP66wj8hObUmUIf0pCktbh4RJYVpCmu9qbploy3A3rH3WF7QCI4TM
/oFwcTC157jIIlLOc2JhZF80euU3Iur8fVcZutrDv9QUelw1yQInffMmg+J5U67+loLSLO/78JoX
4+SKVP8gyJtT7/PUA+y9+n4SFwo9ibEQctqrcRut527zCg82RXBwwE0BmvoBhCG5Uhg3JptfIPMT
N9TP5ZMRzKlZVa3bUiT3dXe1u5exlOUkew+6QGMv1wW/NpbOpm2XVIAO7ziDbabdMEtOOdvVWp77
GOm36yqN2xd2oqkaBYJ95QVCreCFzgqg68Zie9sXWThO53pBnG8XPaSPL9Eqn4oCMxtsdiYWTBmz
Hyogn6NAGtfjwVBKSdESk3Y6g+YR2K8ym9+1fIydJbI4vdkTjXh/UsodcKfYTU2nBI4QU3rXyTOC
WEIXmWiuV4rt4duLAGXLMXzxWytWY+0cbGtgD8lv9+f7PrMZp31XzueMZ1I8OOUe6beiE0rDtwPx
8d8btDQi4DcFnseaR4IhL3iqtIWQlXF6e5jWKR4caJlOdAI/9Hryve73rYY7OGICyglJYnKndui6
mQT/k5Jf1E3hTUoE6eZtNGrlh7WQBQcKoK6X00fV8m0rWPZmYxNUy6FVMnbygxWZAFnKPujcn2l+
WZO1WRGMqf28a7+B4FE1TePTo8IQ+4LkgopE0QOXIi4PeBpV6t19YcgyzY5w7Xx6yDIV7qBNwAoD
J/0+oh+aZMo97/k3aS5iFA70DDn4nmMY16pcRHkHWGlvPUonWreOYg8pAyZnjO/V7+56MCwpcitx
6Sft+6T2ef3MpN2kPmcueKYteX1Xn3d9z8djM0igfPNtHFoS6e7fbVq9LZQuKUrBHd8A8T5WrEcG
MunStJ6wfwOvNlsj7YNGL/7R4R5JjdRdUefAxolcViraj9BWlDSu+AuP1t868nvDa1TH7PkiVYfL
9UwB1WgNeUTRkrCNNgq3EY/NZW8Y15ZpyoZR1WJPqok9M7L2dxLd8yG9bmTfnzVK4gGc+501tOLK
3+rcm8eaL6Pk1mTIakJLT290gNWQt1tVAe0L7XsAwN//GwCwKic6sWHqgaVdDrB7s51ulK6ov192
cu42dSqAPR8VAGjlwMA01FFe2VuvtUPAe6mBsHTox+fTu6NR4jNm/QMLFaLjbX95oa8rXF8ax1MT
5Jms7R3Spva08RoVwlu0KAKMi2XzT5nZjgg5CAr7M7yUN5icq/SQV6BKvLkcRWnT67Wwr9yYD3j9
xISfuoOewNnV5wZHzqAzXcjRM1Cr6wm7jsRUB/+QSwy7wZrH4VMnlSz90XD0nqpPiMPF9bRSHZ2h
dfbSVyK6hL/j7aNQEYzBbCHSvvzsYG70fdeRPpBbwfzpQsgEH465inebiR4DwD94TYqGNBvzOV3Y
mLUQssZllWUgEQkZ3hVKr0VdhbvRXxd7kTHKKqs/ARvfri27GjG1O+tNNCfZxYpMXhDwdC0WLWNI
jUr5XMmOqiseTw2y0/e2niCz4/w1KaZIUNTyqqRoy+8xtjOXlCWe2BECz3LMVRE3xcYJcknn8TkG
9rgIus3jxLR1aK/VtVfDK1PL1e/S8vchINtvt6wmq6V7EzpcO7uMYiGXw8BiILPG5L8FjyMsRdjG
OhxQspzCFbiH4DAn2nIMxbK6jL/obp5GP6Lm6gJA7JSHjUPcUz7iSnaKSIjL6gzvLXQYp7wW2UOC
IeEqtKL9afPUxekLZFCAoGsV96bs6nBteABZkMJMFuuCmweCxOnVl0K1KiOglfoVAjSJOmpXlcoG
8RhbIz1niFYkHNRcgf0dFf0ZWhW6kDGrI+NI9k+faJUUnxloqCR/IWbIsunGgDt6qxltVmzId26e
BsHvBXRWO5bH3dwQI3xPfXqm479+SXG5GuLosErr0qTQX51sBPnZcW8hLGW6n6byzr/r9IK8U8nT
EhFDzNiqqOAgO2OFahf993iBIFk1WhoRH+3FZCpz+l2zgXwysfksDgCXuQJfv4kvpKjRzae4BwBp
2ftOunUNZMDvNqO7aiWucpWpGiuu5Oezm9frAlgY3aLFMbVNxR54lDwhs2ek5OKheIpC4oCM4W6D
M4sCXfMdwO+ILLI1Q1qNlwCWQ1QqGFXH52r4o0M7gQewXq3q08N1J8zZkqo7wywv9O9mTXcubkYE
+eN6lutUfa4p686P4XPhMUY+gq7yNSSEvZjM9VYlrFfxAqSMNtn11DFutw1Exq3RP3RYdDRandk3
6Tw9VnTU3G3fBmle4ZMCk1npxMUcGh26lrgRUUO7ddkLOH37fiBRv0PJueDknuXAT8oYWy5BhxF7
HQQuoaSf0ZS3r41KD1TQpahdqoeV+FcWvpDTpN+goBwFo+Bob6aYiMVxQlYac9dNTjGPXPRhKDfT
Wgy3DwdpvOhkalUBCkuqjyan7hReP+FOuIbTjI9sJCg6bGJ0hU+ocPie+cyFN7udcTsJQaaLnaLx
ASZqoQP+sH4fufzMXBWD9T/6CMakQXgiR7HLENQBCFdUwc0LTiLh9AEXLwgrIBuAsQnrH56yCN1f
KCiNJQCClooD9xwaaXDOnaIz7BUtPiAqCii6p0uM0IyOgpb2NZfHiRToM9GSwbI8Z4e/3VFRJgo5
WydAyuT961fwCDd9H1a21oSnQKHK5eeHjPpH6Nuse1f/OXsG31TYh77ZCkQahakrBMjwSiOQLAV3
0vL+dFtFVGavzyT+v78so3Nyh3X1CwuII1AcjiFy8sGbg2NTlk2Hs0S3y6RXiCdQ4mEcst4PRuPv
gxKI5LygDyBSGDOhWSdfTG2H6NZUbEByIpdX6Q+E7jTZ2/IKM1jMDWA6z/kl0gpREqOdQ0qIk5qv
xgqgN6eu1QCsKb8LQS8I+Tme6mbkG/ZzyRDy0jPj6IWgWn6p6cOOv/YCKKfH4De+Of+PlX/Nk52O
ohsri/wFnokeEza6eCsWtN/s22JOp76FtVCF++thnoMJAokaO9YAnoCttftn2HU5OiX2Jofq9Iig
mrZxu6/f9nuH8U0P1GpBhFpRzVGVo98HvIeSlJ0h4g3gcvIGqWVQ0DSARkrjoHDrR5FF6gr38iCx
TndWVm59Y34Eos1Lah9o2JxPawpnOfpJq8zFwEd1B35ZT0s9m4G5nZC/i2RJDKFWGonPn8pzzPQ9
0/Ug5kcJROfFZXOw5vY7YlXDK+6InAeC6ELspLLZuJLljo2tRBbMxLnckMIByT/preCK2usJX2yg
BH/QyDSUdnoZ5n0cr5kGitlLmB5so5YbNI+16gEN4uYiYTE5PQWJfQYLDnaqY3KuNSya24nbWYup
P0hxtZqh102kkDPPfmZqv97VgetwutEYnx/KL0FC/5GVzgFrU69p0npr5PNCxKpmpsT2fBYz5bvY
XX5n5MranpxnNjPZYdzBeR2scFkK4SgRCAS5KqAWSsljTLdN8LS//vi/fBb3qL0UGLiaZ6qCnJha
gSfRRtRPc2eHFTL0Yyx287wpC3gK4ntVn7UvRIPPULhJeuT58THm7MjBOl0JkiU2qe05OF4bwv7b
Q70JrPPgGz7adTM6qfVr/tOz1xWY2HEQ8Vp8/INuZoIBaG67wjWixZ1IP/BrjyZ8VLFwtBDCEiFi
1TmIaJLVLOT4dej7XTebwka5cviLcXB6hPNPmgXgzSz38WbMKlGFj6/W2dBykFlMig7dR2tOdckj
EPcYUAUO8jfwKmFiDyrxYKwIBLTedguaPtHn2x/0f7BwN+ESNOSpK6+QtTHYEoL7dhAKA+C1a8Am
4MbzlAa2ZuQHWnv27ipoAx0Fswm+kuz2Qb+tlhGZM2TPlDNWsEKhUtywylxkFyYannJ5+ytgwEMl
KySZdvaz7SIT068vbhOZ0ZbP4KuagSVwfnJWroxAfZD7v5/hRPxGBUQsTlG3JiipcFFFNjkT+2kQ
LlDSKnJGf21dhqBV76IM8iBZk948a0KBzpE+fU5sTq9kzL8wgWOe0RZzke1V8qiTCGvXXvSWIp7P
8JJrPRYrPxEifSm29v4zvqO4Y36ss2EtPZO6IMmo4WP6eGZsnG8wJ81HtW4jFjkjGYvXAIWjX0QA
yLeql4Krqk8avsTa+grwhGeCbjAEUWGnHtVGfQvEXFhoBwGPN5bOO9I9zuAu1e9I2ue5mYor9yp8
FG1auHkaACykpqkL/2nmxoXcpmcQApq74R++MRge0dplWb5WPWtmJTNQXLMSe6OYLfbTOZtwh3IF
vMefNb1w6vGeWG1qsF28syqLQzT51rrX8EBMMaMPvGTOGJL9qDWe0b9/FBTfHD8FW2vJ58PR3+jB
EK2NW9O1lV5RYfU1u6tK9Uppk+XuO+6ZLERbHo7FZL4+CgYysHzuiN3XeGRC80b+EPeWMC/G9VdY
6kAXHsS2bDfqNURjdrKKxSFcsv2tSrROtYBrIZphhOkAFi2jcOGuHSpcYYvf5bQF1gziJtbLLUkK
eaMdx9IyZ30V5J5lonvSVOs9PljpqfP63WxV6FURj3L5xYL7MgQFrpmB2A7Je1nSMKITZHtZe4Mx
Zj8ysT+gRpEm1E4vIqGoXu21OEkS3tT4Uf4qYY+2UWzwTc4NgoY7p76OjjdwVT0CtZG1bRMCrLuP
gf+v+CRhTU1Xjc+VPt75sg0YeDiUv75bGxqpWDFVyfVA8j9dtBovsXQntU5whp2GPcKd3aZuQjPd
u5utytY3/loLYUHi8qB9CjalnWn7ZDTkIj6033GN1XFgR9UP5Vbf0NHQMDgkXCKLttIROn+CCqtn
KPbHkVy22b20Msds2EAVg3K46BrZne5JqIOnoyLuFxjC+0ZFheZ6IS6ci3Y3/336+MDkbhYiNljd
2QlcNJNAPCgaVEkGnyrvDMNYyLLf8+dqDxxRkLD460j3U0GQFOFb5KC0/l9yDQQ8UsSq/3ofSWwu
7JNayNSvIkbm4UUfJ2QkVVpWh6/OoBYgTjdgUgqc7Jk+rDeFEYWCc6PVlti1I7qPqKYKQwJsTvQ3
uu2txz30ARYZ7tLdASJfQnNykn+Px1Bmwq0YJIfvtLxxhh2a329w7KupM49a0fd3a7K8ncXSJ3pC
GNMLP/A8KU9ohcLuQ4qVbjvMXkkUSA32rCKZuJS61zst9A2qoRSz0STBCd0+Lmh8dWKRfhsimCQU
nQ1yRQtC/llVM0BvN8FLCqQnZ87GcBsXaHpDUG+TQjfetWysVR4JDR2jbIWHgQfNK3mBq1tLEd5t
SgKHzaXy97KeMn9Z8sp0PaPeReWDNpho+X7+zvKM9SUqtbGtbvBOqyiAXYFnwUdDOo3jw7wapGwA
n+rbQXrGehwKLzcFhM1FL7F08S/RssILncPFxwAmYcm2ZJI8ZuAjMZQ0Fl9t0WCHzSqNPIY94fdW
0g+hUXEfMpALwCFBdyFOmclDrXMiD7wlvrfttCarvFYeOBAGAHr8YCvrafiYMI/gIrEdyhE22xCI
GKJHh7QUdmVKJO5Y1nZm5qb+XhUg9oK0L9TrQ7YY05DOZc8bdErPFC4zYyaYX4vIWhPzTvMGqnAx
BGTfGj57rJ9IB0Jel6xxXypEwB0GUIgRnNsSU46UxmsEhLKUEBxPOFLTXV3BqdDfEFEAJ2yhvwoR
rCry0mU82QUhMH16gyzHRDKlLzMz5XVNq1LbI5gcUuzLNz/8MZks8VEUHVBJ69VUgqfMqvu4wBy/
E4m3mtj3Gl20LQ0T10zjZb36samoxBkHfGVt/j1fLaiZXvb62THGMo8KKCqojEvzgIDOc8dVse48
XdJJPQRwLwixVrQcLR6C+PXj6/Mw8vHNq4DXt5wITdO7tlAAH2UHFdcvKmnt3uE9HOfD8w1nciel
7nkk2J47D6g48WRc7Ww+0qKKi7xvZulfXL0Lm04SekeHWideITOF+tflUZzayuUEsnLmY4NEHujZ
Y2o3bdNL9lPc0qZRtY2erwJw7tLo8hNW+Tk5BOSbTLguPJnR6Tf7Pa7EVA3RNeBwmB21VBrlhdHJ
/Uj5kfvG4/PFNb52LUgoBTQ4+oALKgTndtviLwJ7rkAzr0PsOaQniI3UQWDllcpbHdIX21YmI3Qb
C6suKx9G2s5pkylMTbcbKrrmP3afR4TRDGuMjKSzxH7An4gZJ9zLLilZbcwm/yytRAUZnh7q3Dgh
N56h+o4bi0Q2ISb7aL7kSa6q0qrRmnw8CSL01fvRej3XBJuy5qVG2Fubqcom9pRvOnoFSvvUWqqD
rtOjAAyu0dvyCKAIOKQzfLA401a6JD6aZ6cL36G8WS6xEH6mw9kR9Vu+Loec7lQk4HnHtON6Pykr
lR3cfgEvuqLPTY9yHUb/U69P+aJozo/lHzw+DYsHEa1Ez3TKk0+RGtDnduk9Rtc+HNAp0mEPm7LO
fXuOY49DLWiy46Tca7hXvSresOrHzzeUTLAmzAX0oDmY4+dkJLBPR8UElJ5seiNn+MebQoxiJUSj
5c9Yw378NNzu7kkym90aMLQ1vHUgZDKzOYwTE0ZD/I+xtbCjikFLCGEHyvynU7U0ab1E6q5p6HEH
hNthRV/VE7tSeDbHoQF4vIs4zo6wZpRjbswhUH3+ECshlzA/sKbw/jvXjWv/7h3zkA4+RL2z4t7V
9Qx4uVZT9Ex7vhfx9S8emIaQfWlFNLL+jFoDN+ZmLz7siJ+ywglV2Apm3lKBv5yVp/K+KaSCOI4y
PLkuICIJkAzDEWBPOyoZS1mlg+EwBqwiltLlN2deKrki1DKyOErk16AgScxFggI3ITq2CPkgJ0ea
v2Mpz3XWDYIuJAw/mKKhqc6B/Po2a8szWmOiWmVNgMlI4kQFs63IdUx81k8sigw08hnMHq2ydRTb
iOORVUubtVoNRlfnSW7Mzzqflk6n2IxLIRJHdCS6tE+tb8WNpokJblsOW9ehtQId10D39ulUWEHc
jylFF1lkq36LMkHtqTEViW1aA7teg6G3/ErVYpbJZzHEJbIWv1Du+lDokh6JE6t4LAdW3ucCZtCW
1z3EQHIbUvz6JryaAb3X0gWM/3hkwwrRSiCs/x/6cApYIkWSdvqGt0uOrtyIr+81rKBm5RGBrdzN
ADoS3SZaYXetvPWeEwzhXi3AVvJq54xkOpZJS00yQigmhxRyyAYGEg1+NfYRyOrobif+P4H+qzt0
8jo7K6ftjk+F1ek4quUu/RMf2YnFQoGNJokpKOLW/IPtKJKpZweWTddq7P0S7dAZ7Xu3WDyfqQFR
msS13cR5P/P9JuC/vXLgvPdJleqwVjnaBR/u/oWB/IMU7J81ymIezPOKruQ8TWKWXZr07jMQ+y+R
D86PB6Qdi7eo6xj0NoJfWuS2hE8yt7zeloRXhYp4BfPNzS+AkozhUlvTV5Zg3Rygo0xUDYqlsAHd
snYLH2O5n+XMCKnzdJAILUuZtNzZAxV6sOKuhVEApgdHiumA0adVdXNUNXw2ME6XBXpRVHI8yU4M
IX7L/BrJHUE/sSl5cRv23tUz8q6OkRvKfGHHDzLRAnhl2HZ/PaYqvmcidpD5yVVfatRzecILuCaZ
YyKhuiQJfK0TzGd3v9/tUWqVGtyC9mf01QlKSEpPat0SehtkmtW5wHBrLLj8QDk+LO+tGWWbFHqO
87P58JxMYumWEyYOAWxyJzs9y2DKP5oK8O7VdVpapNVrV8VxTQyo/kP3F4FZWZfln0L08dKT+L7d
GHT2935qPZbp2KeREo2jqAM5GxpIujjz1p8TqwZQLBUTr9E+dCknQf4g27SEuyNWtGV/+9rF6x4Q
OCqu9J6mNlFyX6eoVm7VxfpG/jCKEmFBooTUJv98XGpowlvsy4ytcCfbK0EReB2PvAOX9LzW19+A
NYd8ETctxRXbzCSXJiyiQfaxnvLOkeB1HG0fi5DermW2SYYrhKM8Z+hiHo0ad3TufAy6IO/hXgwz
MwiiPaC5J3VRrNA0X6QUvRjLWUC1YMxMv9jnsg/6v2t3wDeKrwN+xhYpTM6X7cYVMYsfMtnZJMJe
8UvPZNJvmhh5ofbTSca1wxTfFs4nBkJwDS5JHJdI5k86AdRFECVhYNwvSP/fil+jcNVBppMUBSyB
SItctz0X38igeBMLcVDHjid2fE/xcL5Px1vzTopCJMjeLKjvgHrbEfs5lcOcjFEmQrb/dMNysIxe
GDPC0xzPFRzxXSuFU5HhY2JrXZBw4AS5wizq2ZmGNeAt/cZFMT9p6RuIEtZgdmrv6JzbBy7JKalq
1zLcRBD+wQ5gsLOpvsvXAfsOSgg41mbhYD40temRJBs+tj5EFfIVmVnKC6CDREKr3r3E/IyjHeOy
pHEj2VsRnIGv6Xmp4+E71zecsLtWyjMtIxS5jU1QSgx4/HUyV/C+AI2vMGfqu93q/B2nqdOKVQp9
QKPb567EFq6aXRVXKkMOVTqE6OCMMqLCstWoQ/UNOK2MpN6aSJ5myGH9a5+8qnU3pA/N02p9hH+i
ep9cypOl9SxaP+jXQhmDBpafpD/OYyQdWyCGl4/dJm8zQhpZkiFF4DS1w/gXzdPhdw64C+0UCI9b
ePqaES/l0XC8I4mLjLz7BqcdlfjyFRGgtbsOYeHwpGhrNNHZJdZw7PbMT2m2wZciK9b6TRzsabKM
xyTrck985EU1+BWzD49gnQNVjee8WQ7Zr+KIl26vD6SfEoW7ynFZdhlGEfTfevYwb56u9EDE4pHw
6FytKfXMPFUlkCYuBS3JdKdzmIEe1RVvk1yb59gNSw/QvRJh1D2srOnz30qSsZoBjrB5Rmb+d4Pm
Q/ts2Klncqu0VWWFfTVJ42SVkQoRPH52vuIGl02wtkjemv61YUZZmrfU9pQmXM0sjnFgqSvSYQEh
HFfr5RQ6uhrVGSYppAt2bS6Hh+XiJ2C4eA47GTJksrZpRMCb4IZn/JIxLmNjgpmAl7SJB/MZ3Sl6
TQJJXmshtE++b1OfMuDw8LtepgtqmBM4JnXG6nN8O+44/s6tz0eCB6R+VXu4wROIhh9dpCIktnL4
ksWFdb0q29VoxFDiHwUgMiwhBYrXi0/mbfosXHqIfitoXKhJcNwEqAWnZVxhbGfCqn/tuk9HO+tr
5zEfhjy7RflZUuTdligfNDFichiFOFquKET7HIQLsfA63UfAgMizLFt9OH+v7LGIi0GQhX7ecuze
qEUlc/Jcx76Yq012li/4N/y+kk+zus4kkvzIkodohWxd2rpcNznP8LAzYD1CNFs2LgIhEwjyDu7n
xS64F5ATr7xG5abEmnDioeJT4y9MhMEagO9WtuoNlVRgRdsFgugq6H2WT/iRjs0QcuFYmfUaL97d
uLflTpoYU30jPhLEsPgKeGdjPeH5OI6seDyGnw7PY+OL1XYcuNm6icwB22nEThnQzewI76EP9dWX
9KsS9cuaPybbPywbU4Yn+Xrv19CXdrruq0SpjmoJJEeTE3ZcI0vOzvYuT+OBkOsuokTQ3EzPsWhY
7GH50jLTBwkelX08w8QXa9aaWhE5IJn69pq2U17kARwJxJiPXIJYqbh60cbGqcenPS67sCUa+vAw
9J3ktJGZw2YmDeQsASsRs7M2OcWxC17PiWvwyhAEQZ2p+Kl1sd1H6SkVgfOozbSlzWQ3x8Uaqeds
RRTW5+b9sDyUIUFeXr7A7HhTFZg2kvJThXACgNxKvxzShN3fyibY+VyBiO7WBi1yLcU+7566NsKp
uMj/o6Wxsib8HrcraPBMPvmMtQG2cvTFOv7P9ZU8FEbf+UCKlIYKcOKO35lNsClmxw4ld1bZqobl
afb9AY6LuSbVH94EDLlSCmtFxTLgr8eNA7FUCEZNCCawKUElS2jGJrFbJ5mpT04OtAK7vi0NqyT6
3C8cElOHrKyNMViV01+gusgNZoCtKwWWP3kkagqMWksC6gBIVzV5XyqIGXYUFzTC4q0WQ7Wejrqb
wgvnpCOwMZuW/fVtnqlfAxSXIo/bTbYwo0bzQ7nAvauU6YdwJjhaN1TEEaC9cgiWbyKKzmImuvOS
o8uKQjnf0FVxEBixZF1FxiTZeZfPJ3sLfyM9QA2JbY8o+o/ruHmpalPDQ6686LAeR7HrtzsyQxwn
/NVu9T8w7lNNzWRcPxLIm8kJp2q4mQV6YRmZK0gtLtgxh/CrWF7iLX1qF1Izkll2uF1qfIYoV7xN
Jr+Ecc/HRydayl4x0tzcZ9YVc/wWAfCR06HF/9dkufjaAb/lP2T/vX1Bi4zYNhfjvP7XqPyqFaD+
8TOWsf3FgwzseO+2EUEMD5z+FmTXAggUNU3HNrtMLV04q9hHypyg6f2lB4sGAdtfDRCmPm7KOQeM
YC527QTVqmUq0kAYr00xThCBfVCwDkFHHUVXfVOjZxgUeHlOoNGkPLtlbZulA9oG37DuY6QwGtMF
ZxL5Xf0oQhoPKPR967UbdQoWiwWlCpmvW0WtBhWKvUe+R9J1RQwHThu2wkaVXo5WHsANnOfXi3i4
W7ievvHakMgf4/9qKAA8LBrks5Vaj0fuJxol+fRooZ4HHSpsCj/7CvqlArZhEBKNZ6KWAGYRpR1j
EvDNNvMpU025PiUPEzr2IQXgkq9TqeL1eKgK+67Aa14nf+ZXdAmiBCwUXzopqXAldx+FUG97hQrN
lokFqWyHrtBClhSzodrWGMwzk/gkmo1sHevXCouJg14iIOXo1Z57Jl9xyKkk27GwZIwAIfeBe07O
jPhfvi7d/KqLBbbDCAV/6NSoW370QwQHOXbziB/g6tYKGJHDmQ8ERZGS3EvN4mQLC/QHYoxejbZp
/qkkZQgreCkXVuJ/jLd9xMVxMJ9KCyixvMLwgOLTJX8skO0WVQ+u2Vl+mI7XlIfDcv/Q7W9s8bXY
kVt1Byo6KosJ/E9UrTEK4cTbETRPZBEaZ2HZ2GYkWLg/6Sxh7ts5+1K9qQ/RuvYyiGNuUyejJnhN
WLl368nMCpRHj93SqCMcNo98NnximaudRq4IljnuLAe5kRI1izx9kxWA10x1KYX5xA1QVbMu9WqD
qe6AUSzVZ1aRa5CAfYnzInBOtbYUjM4AV1MOP4aXgIta9Op06cyo8eixMirGRO/LeWqOlFQFei2k
ttjywjPLnTZc1SMU4yhSrQoN12xExYffDeCShMt64OHvM8rFNuIxoe7uTtYPIqZFNnOoF+/O+xa4
w09MRK7Lj1jTHeKfF/+xFE79tty0tNizKGFTIQuGJf7Hc0zNaqgmbAy3EntRZ4tjbStNFf9lwcrF
ahuGR8L9AWM0sfoGQlB3o4vUHn2Tb3nPC8wmwkGwR+5zMakeWOY9rGeYVpn3vFIO6OmokZon1yAt
bpDaP3sR4XrL2KeFEg/ckMTTC+pS6pMEGVaJZqmpUERQnO3yK/G647il13FqRBPkNdqMl1iOeFCo
tXcsusek4Je36KiJb6MMh1AAB6SlSKHAFMGCP2JI65RnYf5AKULZ8krhewnM421MOy0Lozu+NPTB
Dilz5wSrXk7Pyw4C9igfAfL+DZOkRPUah3D1RChgxQLiL6Kyxmyasn2C3IDMIrE6xlpBDZ5FNjkO
n77oaeRiOrj2VluUtvEstyIicx95WpufTby/gHL+RXsoxqfGNBw8XbxF1u+dnfyLiuXzBCFKe/AW
zCGbX245oCRz/FK6TKSfZJJLjHZ6SFI+ZItY8izSUTapw+wAVqnwHbeDLZEkxitGh6SpMzsrvyDN
dcUTGVgzBjBwLF8TNkd+izUbM+ZlsVPkZKi1dFRvr1y27M1XduUVejFLAd++XEyU+hpK54ZG1hGO
IkSLbKLFRjimy8nUgSJRb5y3Lg+rexNoFKv61a2xMKnFahauYfyLN0xaDalK72yPa5oInr9Ctgpu
edMFIa/4hMPviO+Vu3IiJ3pfyvCiWxb0hf/GHojMskKJQyRyME5GtokPX4S/4NxdWZ92bGFVw6z2
v1j+YlGnITabHBjdNXneVnbd0qxbF8vWxNlks4Nkef92yEHvZRQqihlNbubC1Hz5Ifj4/mEJCORS
vnN9ZmjN3YQznPo+9P2bPzZYoKlkkMyDmrpXWaFuDTeG4UYaFoxET8k2Flf9Dom9nvpE2/zjxqGy
p2oouw0IoxtsZxYeg0/Rkl86DMWWqRMohZ50J2RKFyf7X0OaS3V9mH4ZEbE3H2wKJyMLvq9dtaUR
eb+zpxS3UkqhKXcF9u2exygwso1TdpYcPQBcVKrjy6EktjKfQG1AMK6wnMgExVIk5O/ujNhrhNDT
ST4vgSsvgXhlOWRNkRjmCWFzXJ5A47QEelCyHuAcAcuqXUjNAHbtQq215wlJBtN2EVf/jpORsHzb
UnNNJGM1nwYps6baCuihQ3xnbqAIOwJwAzCdBY2sHWgW0xbfwoecXk4PVdjmlyrgJ99zz4h35gEm
r4BeCafYKnoOgFWC8VomDpbQFZSyUDGs6bDe8osNgOv+0KLai0Ys7ssNh6eTjljtHKOXBtOZG4sn
c710hJvqgE1s/DaQqBfdDS6x7VRSi86cQYs9KdNMNtJxpsk0CrYa7NSBTr2lxYlT0NOzvoEXMabM
0yC0mDv4Yqk01IN3Fawnh1WPwumURPrs6Oi/zsj52MdblDhVjZgJEtAHIPQP7uCynXC722hmYud3
b8FAUA+p2CvztMIOBNFDIIroXI2PSkpDRg6hVND/HckoYobOhDxNCvDLC9VvQUBzW5osW90zfy9a
1FjOU82Aa09TAE2IGIhwUa7RfMaE3u7nlsKnHSOVYkR6Gw54uh5gdngFmNwIBzIlrNfIWxOzFRn4
YEq7a1UuAHgN/x27Fu5vYdh8U7dd+A1hkAH3AmmGbwkfa0mcnE0j/5pMhEV1K3b9GLe+NVbpQQe7
Z3gsSJqx1FWC0jRoX5ag23xIBp0J0Ff3MygkSmvGy5Mn6BX80hzFippOUH5LdkuCiKC2J5Fg93EH
Xne+RlQzocbkAcAD8mdKmbr+k06i0mm6QH6VVXDDjU23s6h61bNgpmwV4M7SOwNfuChrlRS+9TE6
ylSQIV5leAjY1epGJ7MqEGdnFKa9PbJ4kh+gJ2+sl/Ira0cFlK1ZaicMuqwPmcBd4upCMxizSlJC
F1ASK6S/bqZKFt2sEE1sgzb/hbBPelUOykH+UNPqYR6kRgF2SyKUR847js2CYbL9LqctbKSaLDVj
2ICna0eZneZq1NszFL/jGDNszAycbivecjPWtYFDlXq7oJW7L95cPFEJ7lZtjNr/Z2QsY176W4j0
u3WdzGRKIiFJOOCMTEo3kYzi0KbuLBfdy+yObq425Cqx9FTOeZNuww9wx/BEKqENDc/E0m9B34Zs
B9482tcEIwyYc0DCtPG/Yzl4bwq9IU0DSrZvoZqnCnnaVpc+6ed1b9XxvjpWsS8plDb6MmGAKrAe
Zx/X5OIqCDAxgYHCjA1UmdtRwl/Pi5R+zOJYo/3jywFvwt3hLScpKPujYZEzGfWQzVOIFnPnZqO6
faR/x47Nhj52os6VAXrjgnRbIjtudkYgLxHnuEFWM7dTODZv5xGtAjwpqT7b5SUHJB+zpjCgvcx5
UVywZMxhWclfQ05rZIvOlqfN8ekZVRBryTsRo3Fjjca96g5YJDBghnAt5h4iI31n50X6jgaNMDTi
sN06s/duTIT3kCHhnJvQtDln/+Jm7yj2AuCBYsyuPGocoMc9DgSjzAdXNn1+vr5lnE5CEySzTx7b
PAyhM4d6r0sBLSqNI1rRcmxdFyL7CJGk+wh6FIxJRYO2BFoQ74ig46ygZOgvEXTJkCbYNEohi0i5
v5a2pcNxhfC+xniYbh/g+A3QINzoqkWDWXoI73rEcGx973Rv3lFgFp5oS97Kr0AXKBN8GlwvmMDK
YSYf77rES8iH0j+yk12H6A7/gszVMxyoJlYi5gzMQpNL4jwUaSflXWdZK/pxLnOlklK/nfpFwG6z
0s9VJ8hMJqvvc9vbUhk51Ybtcg8zvn4Glq1ilw9nVvhJTzYXTlndCjVuemEkq07Lk6IJNG83Ejyb
GQFgfq93FtZlF7edvfin+to4GuW0zg496SaqSoGzEWvELFGCz5ffkbwruoDT8icC+fPWspiCdjNH
lHS9f5GaA+AwrgMIV37e5Zg2SVtdQFfblkpdo4Y8cPP/NUNSYcdeYPe9st0kwDqD995c1aPwaE5U
v0r3QI8tiMDUh4fe4Ul8CFJx3ZYPUEr9sq8yV23w80ty8gGpT/508IFTBug/mzedieZjk6t5pT26
dN3z51KhgKLLnPqcxLJ9Vtm87p6f+1HZ5aFycPz1IhHMtkJN49ZR3szEEoEiwufLLyMpa3t1weOG
Tj8ja7nj8BIhPHUz23ZNuETaX9PPPsKeBdaK9ZzW0u8AOgCaerN9ob0vZrE3EbR65Tep4gHQkhDX
azDLdUy3ovJJ338ng9ZjtuiykuZzOwtUQ8WRhN+0MY7+mgK0MMaZ0krDceiBDgS6b3Xupblv22sX
yxJSU+ukw9ksNkZ08ElLlq5Bbap1Hh7Imr6XQq1pgNrLJm7G8kh+0lpb2iScdKQbpTwG6r17cRQq
mumhyLNuEj1LhfuU2urSppNtEsCos3vHqjBDtxI6xRlv6DR79NlF5QQrtxuIwsTUG0a8N0WaAEVw
yNyWZO3CWR7LqoayK3oejR3ssPAW/7nsCVmCkAiIzhKAqMLLTHLm94+gBCfAswi6DiViOi2vH8kb
72AQ+YGZNDjnKU7YdjX7gtt3RWHt9NGHIn3+uaFeqmHgRwLEetUiLgOj5MY1aRr9VYTA4HgjaciK
byJjvmT0W10sPWVXNp2J/rhsg8lc370HHXvWu0chBkZP0v06FWbLd6lXFS8xZb9KaHeQ+PBN1Dtq
iLlBUrjKpUxBZKSPme8kxvTCwdLMoOx7u39h2Jn3CcsTE0quMEuKSi7ZMPQbpi1XPXFe3I4DwVOG
gPPm0K87qg2kehq63sDgdWTaudcE7iiOfAgXKR9B44aKSrZI0LV6VChXrYU6ES8PJnNDuUQpwc43
pXrlevJioLkownU0OMgS24/eEKOx07kYus3buEIlMKx3PyKtZFE5IiKrsJE1Xh93WnL0RUuidsDo
vY++NBqxrJhMhVmuwaw4MgpxY5S0vtZS0KkvM9A8mT5KGLqHGsR0OUTsYy6/q09RYBw2MD70iRjy
1naLT5/l2SLjZGPar6KHwW/8RxD+yB0HMPeTuygUTmgypL5Y1ZMB7dsJrN/UOArjX11NZlviOsdu
5zgaVsBapn+xWt9lbLukp4/X/T1jiJ8Tss0J2LMV22A0I9mrWjuRrpsTve51o9ts2VtndCZgr5kb
u2wRfGDWGtkjmo/ZMf1KcJw22E8e2bIPnRJoUmuMzkTKKi1gstF+n7WOThcCAF+hJqKzgbg43tzE
tApvAJMRBZ67tLKBzUv8eiPEAh0En6NJUzJagqHtEL3diXlVKikKz8CyR1US6wDqpS6Cyp9jW6/N
7jfDIh+ctOk4gykKufNZwoEnjWjoeNrR5jH1EH0uf7j9VwYxHA5x4FMoXZDcqBpPhwPBwbT7ubFU
IAS+LOzObMdjdgGI0nUg+Db/RIY02Nh4w3zKsDiaJklEZWsJ5vRggb/mczbs6C+H7/xhM3xQBj+n
sQEpXei5n55usRZ5W0EuUDVrcysYDZZBm90a1xil8/yMxSmXH5uLQA6O5Xi+g/8qz/zMNtQH62Oz
F+SP1VYrIC2fBEVzuRm2KSeo6DPMIiVm7jE5w+FHwUe2LIeI60Wz5GixkFWw/HPxcvD/u4tRCrDi
9Cs9XwWBSUyY/XDF5vDntgwTrwKQmeSUZNSOVIMz6IQ0vPuHdy1oClPHU9o8XnO/T0/TkXUO+/6F
tw1j1WWdtRXCEnR+kEqi5VQrcNP670Qosv3Cdd64wRo/Eux3ZgoykC2I+59gLNsWyr1hJDQeXScV
kBmN/dZGCdUJDL969Y090/fYd+2JtyJYVsmAP63dgV3kUzZoPnuqR7Da0dvVB3RSld5e+2ejl5Cv
8HeS9xY0U+ZkLQH+Lkn6jd+k10QWoEN0gauabzZAtDpEJDtfDKhYrtyI5fFvuc3euwH+0qZaFzEm
U4PoPqRC+m4nokgp4L98Tbvms71oq1XVpjlCslSmk14jcxH9pLY6b8/dJhVZ4gIm9N6pTXLVxdZq
5Qpx4ogN+9WPEHc9Sq2+3J/1a9/8s694LN4YcJyibcwGvXjpPT8CTKTAkpxN4O3q9yy2WC1JMMje
bfKY4hY3MVREm6xLbuUvKgQVAFXXYHvQ8vXIu7JMCeLcIhZmgtxbpzbWA7w4touukxrCojjpN7eJ
Os2s74y4SGEvZHhkBg/2MyTp28NKSCbwEqKYUbXugcnzNtB4Fjj/M487jr5dO+fJNgX3dVb3Kuy4
ZdFOwvrDt/PfnXjbrH05SDTj/HgMRmk/kzRFoG2xc0sjBnDBjLJ0RzLyq6T8aJ5gBrShyJtCeRQU
L6//oJ/7MtrUeamLYMgyEHR0e8xaTv1Pt+/Oi1wUb6QbPBjyXzQU2UL/6pdqDB/wJtDgcEIErKcp
k/oewTzePXuVSBM1VddhlFLj9HjZ5TGAtm+Givmjef/90fitnbEZ9Y4ayxxeQvSpjRNF97AXGF5f
KiP3QrYIl6/JZEiiDC/M3D8KhXSPMIxOi6iHzfeLW5F+OeAesr9tVPSCrjEyf1mmCQfHbdqL58Hh
qnWSPc52AAHAqBglvcqrolasfIymiYhnQzb6S0JictQ6DT2kj+4d/S8n71w/P+FtQnZ4Xth2xmRm
akh/+FeBl9ANtaShUrh/UtmI/xTxaP9TO5z/S3Y+Jmg3uvhV5S6aWlTVC9QxvWU3c64lw+CaCAVD
VjNfM1r0UJFhseSuoBodheYm5SdWRevJqpzsnxFsvy+M8YnbxChJT6C5sMbMQ9aeac8eDx19MSg3
5tMDbX0i+8zQbkqVeERCIgA20K0Z4yIv7AxzqlaJXFz7wHaXw6Ig+bHLi056LAwCo2xJAp80mwO/
qcEGD8/zhvpl8wwBlwdnykqdLnjHS1rqt5UJvIJt2EODDm2I4Ri+YUV+UyMnMhgEB/y8yQHatHxr
6etJk61iNFh2gjttQv2kxy0toqFfkLEbJmwxuDV0Iwx/3/UvPgZLI+/ShHKn4vUIjLSlQghpOoqr
7ScTeY9CS0Dsilb8F5c9xwh3aYIFQDvohf42VIr62qmk1rO5l/vnDALFe9x30u8EExF85sWe2nsY
u6iiRS6WTiYDuVcJsPwyFTjLHUkAA/DjuGW4ULepsIxbIZlrxm12/HrURzsyLGTwzCml6807QiSg
rCSHPWwiVMCKhi99MLPGbliRW7QF7GDJXefEtQdL6On7oTm6Ihy8M8641rN4RmPvx+3SbXoWYp3d
Y6z/fy+N28y4XDEYchyTCZ+pdQOU0PZBA4qtBL5JNkWeGU05A+EoCWd0Csu11BbpdU1CK5KPjDcm
s+JCWffF09OqS/VU7HxgQEReJLX4N+XOgrvxojXmVLyU1da6w3Zw20BQwPdCpGzBn8JZPMTNMd6r
VR2bNukh9+uvVLNs9LY++BowGX9ckLh7k0Cri/k4FfobDJdrgRsWS1LPKpeKWwdDeAeOFMEUu6iZ
4gU26WOcRydmPUNyv304KHvn9TXazBVN1F8I0VHxzn9hUPJSB7D+YKyks/MSM7Ix5w4f5QKXIL4e
O7oLGETA71RXfi6CbuywwGyV7FW6mBkILjUwlkyuOo8zYXinoSoBqDx9aMsGnn4VX9YKZuC0nzj8
yc/vYCF/75Kes2L0nap4OQljLTKfKc4art5JAJcw4HSD6QgRy0j8duptWNHyO0Tsvw2WEr1kIZAX
KAp6ygg5SFN9ZaY4b1tsg5KasyskpfiPHSgvO+Txyhdwtk3CT2FeywPMC+L9dp27c46eAiFcmhu+
r32sXb3Fxvvo0JhJ0P7+fz2YchKa+S0KEi2vZavf2A/qF/GPie8VMiSSQbdfelv4nUINVQWY2kY4
D3oWtGhuZFggp4DP3BJfuypXKNoW4co2Bwufpmqqn0/2Pb47BfwBJTy5Y56YcdEn4BvYWTzPYZ5B
TiNlPwxmPRfzPxzS4qLMINIAGfUHRKicGIdqvaJ9DmKsLjBOl427hpm0ip8HlMPIKpW2DDl/MBSo
wsqeusZDCh2hqcYh6mvImdDITPFT5iMaXr7Rp0Ar0ANWUQ2ejjYgV43JEb+DAF0rX7I+MnEIwnH3
O8OhR8PNUMDDH4BzN4GfouXRYyN/Q90YVx9reR9qHfx0XWntoThiWxxYni1oePtvKb1V3Voz7nEN
csz9vBqlwz+XevBEAukvIM018Tjsq6ELicC7U3bZLc9cK72I8e2CIJsbAkr9XXKE1uAyDxdc0mWJ
d1x8rQ64+OgHAJoWz2NVm2TM/Iozwx1XIx1r6tJncaks/98bF6dFM4dO2Dg22JculIWy74wr5XS6
NaD/v+/VqaJbKVzYQXTJR4GVhE1jZI4aq8HA1txl6Bq5nVuQ++DKfCOzNnnHBUjICbDzwJXCYbBO
uGUyGH1bdAjYPVzvbU+nZF3fqkceoWDy0GFz3j8G7RjHIT5EnAWRrf5+QnM+2RKLMF5BbWge4JWY
mTQ6ks8ipzCo1HCLKCfYtfyApNM7X1Sc5K/tliOAs4nEMzGan3tm63fwo4RJR1SDfKAR35aX9waZ
gzaU4Mc6CmCX5nZvz/EERI7U/aLEPwwEJahKJbuYJf8jau8UD+yS9E4ntsNUFU49qX67paP7tX9A
uSv7ksc1wqHcFMCkcgZaIyqMjXhlxhljxr0yGWczyfLtzhu32fj/6wDKIvAbubEZnGaOojtqXqg5
MFWbzQrXzXi2eIhVOeTtlM04C48xJOZYpO1+XXudKZMXJ3IduJPAUBP+DqXUjVdTq5dvDqlTwBs5
ecHZx5Ba6GORz07X0SV26L1gehf3wL10aZ5fSeNCAq5phYvk4fM7H4+LcQfTrQk7EwBQok/WuHQH
6TuEjaljBV8bmAIYedgRPdytbgtXFXRP0S3yXrvG4AzJ+5lnqeOo+uHmY+QFexWUycUsGztJy2Q4
21M+M8iM65jh1Agex1H2BDEbBBqN1CNCGt0cVGDkrjOntThyXWzzFZW86Ai8Iy5DLvlXE1PLjjN+
0aIFhfrnKR1ekbFn/5dh8bjU1U2EAlO5NhHPVLAnBYKVqRuSyAPDWkbzp2qsbrWTRjczleho/QYH
lNN1gcWNTNTG6b86hktYcJvn+FtC4bEDPhIM2/v1KTRXqPuUfa+lSLxavAilOuT0FP4l0Pqd1SmR
E4p6zQ26ShBAyEyWahYXKPNTVgqNLIur+/CJqGNyjyEzveYvlVHPqVXbKD9yzFwLixYNxj/q7Cfe
6eTIVbmnSSyVEziYZq5RZ7i0MxBgeTWT4ByJ/UPjIJxEsjT1UStORLskq0RtJ32SrsgAEOUeg90t
U0FfLSYbY2o7392LTprisvOBRShv2gvZSj2XnBxQkEU96iZ7+fudr5qECHKBGVlvlV6Ec6OEmrBP
EmO+rXfh9dG/u3ZQTeOIB51YyeVXco88oFumU1UnMhiXT4HIdiegkeRqFo+0pvChCQ8+U3deHlBC
YvZi0MKMzsVFR70bgVxGyzsg4h7nZr3yz7dlETiVAnM623gRzA5dSGOTYDBV6nMK444N++iN7hd/
MnnaDDYefnrAxUxj2UioD7Cw5T+k6pQX3RUnORhW4zYSSNaAqm9WBNp6xqehGaFggifhuToV4W1t
TjF/Xj1OZof83QYNukdBHTGyMRYL2Lf6vSXbiSuukkfIeg2XV7wsB+Sy8SQUsnbzp9IPfCNB6XjF
Q2uxkP99q+eQo33NbD3iFvvQ4mKuFsfqdYsJWHbuWv3CIE1wu1rzXa/byAkF4saThNDjAa/n2Ow1
LpHWhknVp8/0+yNU0rbWiEtirgS1Z+Sl43u8wvKrUMx/cDp+0MJ9/D3apwWqppE7I4cD1cW4dgEd
OJPmKSpzIPaYpg28nQdPDUQmPpO5xqRgU07mWUFXOAZY7CimGtd7XQzWB5UyR54gPOw7Oc29ub/L
3IYb5ovljgYE+F7o8VDPcWo8sUS9zAUKZ30Aft93npN9obCUK+QAQGH/E7Q2kzmA8l/XSGsWTS3R
CWS85OXSF/IB7Ggryfbf1hw4hnjZTcuDessRDQuMoJ1jvb78nkWFhjaB2H3rqXErsDVLQCaXLaOS
5TTzfmM96E9f1SDO9VBMB1DVov+qR3EavT+lPzIUadY9zsA0Xjr6qGRoamyES5nBtOTeZKK2Dke4
fR/0Ej1lOjKG1uYmdrYQ8tVszo0XZtOKTl+b4l3Yj4mOGBnvY6V3v5ASeZm/81RqN7gXz9SE+RDW
eIne/2gFdkDH/a2inbQeL++KCminxnViqRx8qpSFAgHNN4E58titM9FdJ8fQK1K8mH0SJh4efsgX
KzA2TA2QSt/ialOp8UueWtyP4XA8IevcpXgfdiNY5XuOOSPixMJnWX+T/ZmVMFQ/QibRlc7x4+Mz
mfxgViXY62Fl10+uOu09fg/8fOh/+iOKW0mA4azE0IhdQkR3TNrZC7xS6gLTwdlzYmSOqXibfjWk
7fBSTg/o7niGvaJEF48R4qKxwUOqyEFRYYcRu5QACu5qjSYEY7As1a71nLdcDjyR0Y+GLss7QqA+
jJzpDGy84qBUW/MRPAO5ne5crkgmQ3bMq9UirYtE5AkR6lKzkcwsQdKe8WMG3JH3lnjKfc73wFxS
7TET/XMmDVfXGc6I1C2jjp4LMPeTLqxg7rveXxclSXy1lUBkLXJeccegKVpWKOEaAzjjoJO4UN08
hW9GyW1AaCPthAOwT1Xdm/n5MwhGl8hRn6v6PEeggNmIyamFJMBLrtblV/6+4dR6gCtEO7xHC5fO
ne6OQNaN3x5tTexVMg7k6uKSe/draCXutrrPQlClD9VWu/afW/nFV9DvOZFAzRoFZEK76OORf68o
K+xrWMgGn+Yqe8I+d/8ApcofkfRkt1sWQl3iffDhTj+2b7Sefx9+UjESe/L8HysfP45N/9DRLldB
yllSs89EvVYZWYNp2dPqd19Uf1/Y+vIrAiKJmsrOjnGMr4W4HmFI12KW1uJPRRChCaW8g6aYTGb7
b2GkwK7L8pyyWfVO3DitRaew8UmoYHQiOiCSeWqDf7d6Jjksh+sLoHuxupH+TRRU4vL8b918si/p
J0Y6hiyeM3GvYcKClXHAdQPG85agS8aJr0cY1cmAs4RMZruQaaHLS+BnsQG/a4F2upt3mNE+Y4Gh
L3PE8MVnqlqoNI6H0rxrvCa4p52PTRG4tyf8Ur3umHYZtJEmHhe3AacNOVPUsTn6tj07QGwB9eUr
m+TIIYZh7yiMgjv5b+pDF5ZCmjijbq/PF6zy+T046l7ywzWgUEVgW91bujDZWWd9pQ/ob4fIv/B7
XRIwCvkUoxpD47skD0IqUe+8v2IbAB8S3vB7oS9Xr0c0Ywstu7APHpiwdoFp++m1lolR2nfU2BFo
f9B4qdOD7LtIF5OSMp2/beDLcVd9Ahh9cObZKNje+XaDuhpimC5/e5wrruzSjYhUcyZ8KgOXjfIp
cbYUygcx187ZSJst8Cl+aoORK6GS8YjITpFm/X7Vr70STZ3MrV1EY7SzcZ5X5KCZm8SGplWDAM/j
x6/yCoFPRtPvWPZ52YwVDUg1uu7C4JcDazsFpA/fFRkE8XezUtDKF2jcXyiTDG2yjScTnqBwfpZE
q4UdQQ6vFi7WzVV1KMrosx5mb9d+CUa9KjtCgxUhMIEK8RxljBSYvRfOHwy9O1OtT5IlSSDGj3Fv
vUfKv9YxXXmAPq65OvOdAbjn6ccnhCd/cEeAf2EvP7slm0PLKVY+btog9lPU3ecUeQ6aBKDpDM6r
69dIaPiZl8o9oqbGzutrJAw+MgiXot4AETmtgqnvV5pT4FfLiLZneMe/j2lbACk+GD2cSFoU+jjQ
KvIojzSHJJ4ckZTmZzUdrSH2ak6+tNiVtvONZ69TZ7KIbj7tO9nbCL/li+AfLhroHRuWGdj2QRSh
wJkfWrSM7Eno6KTGmdjLmkPA6os6cCtuAxiCWG+3ZE1kBUIC6CyqetWeWPOHUmOlioCtSDppX9fl
asW/N52mMBwb/cSU6y1yOtCx88njNRQykOdBuQERVjwSj1Lk+0PmtKRLb7+KGLRUPnXyXjx3+L19
tOu1XKvBYS/RtnX+TRveLJyT4KKvAFhX0sTPkyjiQcZAp4jzHalwhpOX1V6Bn2HUeMaQnzekbBCT
aNB2o8FspUKhkTH8l/N8UV/HmZ95L93eqKHJFqsX9teMl1XTyijNP1iZa/bDf/D8UOYn56u7gwrt
7k75pweJNQqmqBGr+d7FNL5BA2rJg4MGxOMni5yxkoFsUNPqb5KJPcGGxhapef7ueKmTvqioMNp6
JtQcDldI7tRzRcQEtEf8z5libS4OHk3z8a9bsW7emeCoGjuhybaGbI5QlTWhkKAS+s44bw8Xl3YZ
0AG4YFvRmbSSn0j/UFX8NVh/5wXIuFnEBbyGQyVWHnBT4TWy1VAcm+PN5wiwhQ+GX0KdI6kzyI7/
2rk4A3t33VQ3Iatdo9TUPGdrz/Z6JppuAY3vpKy0HWgPX7UYQXHcL+ZeKx7GtWE+efZJ27jGniIJ
t0ybl8eO5x0pOObi7Npbm/IzMHGDC5XbZcxfupVV4UJ/f+CdushiBntiDaAurp91O0sq/6fTy16y
uWelgvuVhsC4/EGpn8jfuaU8T97u89h7wJGfeQJ9crVVMCiDWAcNqQRFrZP9be+sJvfiLNoj9Pu2
Kb4R52sh4efdouHSdbHQ5oHD7R00Y3UVvqOs92idYKFm6FUXw2/zLcv1gkFAuMITSzVUMclP2zgX
JjdhwvmlUolYAgiDjAqajsjivXHM6rcTDmoDloiPP3dnrzeMXZ/G9BjWoDMaFrfW5dBZSOM6vSVw
YBszZJ+ClAEcvR7rOX9yYfedxvrsciO1emcxyfK9UdY5Yd2s1YxdCsXF1lL+UF38gN/ASwCyfCbx
pMw8HCXtbRCgc09HK7AdGYLuW6o/JXcYexFypnHRAUzxNGHuamMfduZRfd1aNuPN4i42hFiDgizm
aYctAuGrgAIvHKqmIXk7ZTHHldA9gDL/3wSG/SzrCD6CogBPIoZVQIVhefQOa0/bQNB/zaQ9LA/y
59MZEuv9NY6Sok4cM/Ui9dKdLw7AIyAEbAjdw3BKKBljWZV/Y67rM7XpebSJyXs7nqMLBvJkflzW
gmwpuNJr5h/pAWQGgwYKvq/0ab990leCYgl2GZewnS22S2N5VFGz6ZAK/3UCHJCxIGn2ynI2QTfN
/k4cVaAlr+dCPr0MU4/4kiD9dcuZbaxq3ozq0fXvQYlNvUXFsPm/KL96S89zztG7SGdVCuKuPg02
mg0p5Xas/5quoaWOyh+bHKfFDODzeAjSFvyulGwrkWJ5dCQu9sF9V3xQEB4fmHa/7skteCWWTzWu
jfqGBRw6BeJS3I1n80vdRzMWfCrfviUgDkpbhUDVd/4775eVc/WJojrfKKHmLj74Mpw5DA6aBjXt
Ya1/3wndYUBvCAZtjdT/iaxbDsgPsiLNA6Qnara/Rjj8VhsqLP3t/vymetBGXh6EbvqgP4+k4Tq3
v5KMBC91TUcUNV1xXaWpaTuUqeVnDqIKblSkoRGAnG2ZWksYycEK302f4cK6Mb5onxPp7myr6a7g
Q3fc+TT7nIuKHIdgn+a64e6ybv6lnwIURIyUH09PQvCF3Ofo6d4QLYOMhVTEBsURf8RdxpKkxEEk
+HtAaZbPxRI3Xdil0ucnC2oDCEOg0Tj8LJB/bUZCy0r04eKfWveIMyU726H6jT/g8pK/nI58Tj0d
gaegrCNUX+Oj9q47rx0Hvr6FQR57XLJuEj4pWF/6iQ9kzAhcsbrF2DfZVmqFjENeq1qoDnaDf4tz
pcz8R46+Su3/y23iq3E2rkM2bs0rUpsFslI1dbmAj4y+lQDfdzX3XWCiorClgVMx4lhZD4ABHfF9
sIHOqt4f+vAD/5vWBxRWVmihpqX/Edz6aJUPQCw2yafNHczmnKEx/zqWKfOvtUHnGHWpUNVoV9cy
rQuy9HghiuLfJLVFkoQP3B97lDVghzG+gff+MSWk2pG9EPQiWNB/YKK+GDU+zZLztPli3XZB4dh6
JJHJthY9+UXpizne/yeR0VBvkpYX5TgXlUicOEE+ePDr7Pv9ehDAzR/F+xeNJ6BuM+zJ+NlxI6eX
Kuig9tVSKWWA+NDGZqEck/8QbGqKmrRfEx8grU8P+JWzgw2edqeVfPvgtXPPzlNhp3XwcS8Kiiii
++EsOMxkXVHH3Coe26M2La6TSsuRqmWP667IYYy1hI4+vVRfRZAf+X8xBxkEoKqThQkbKXv79RTT
PTaEor9rvdjqWklfFLgPAAp8pFgS57AgDC5D3RhBTWZtbNY0X7Ut/P6zCcp2zkOC63C55S8oE2Zj
JsygHMu5fBDrX5UO1j1JJBYaYup38CXJjXohPI36RZ+KDvi0FIHEq9rwJkfBAr1qIS4OJ6EQsXj3
+Ia1yATUuMQVprUd+s/axCQ9KmkxkX6QxEO5CGlLGx/OuTv1/YecCv5xyQ4g/LHkAOuu6xzVcEJA
JWoDhCYGlr3jaubWATgqJkCFmDsIo57pQF2KkVdYsbkyHYGoRi1T6TQM9AlFpHIypLrbvw8+3By/
V0OGjGh8tgrs+WykMPa07VkGZjZ+GBnZxp9Y72KnKveaOLdZe8mlLhKwv/roXXKre1bLutIqLed7
ArleIzL7d2lt+B4iKckT4pEMjaKPP/VXwwUGCotqQczIU5z4Kf8le6Q+D86F2nC339wcbI/ODMRp
Qp5sfFOPBjeFgXuRx8d5GuFzs+t4jWnQ1sahKKpjah8J67hNnaFyuFbjpL6GgJ+0LKDjZffrSiW8
ZzCi3vwCsDT/TtQPvXwYVa3Td0aBqgVPM5U8oU7O9oCId+JUrd7F6HANtDNYxcMT8pTzWKKofh97
Myo6NSnKvHfMJ1JQ6y+DkmO18f3+I+bgNNMCvo0KpHCzj4SU+o19bCA+ae6lvu6IO3kBNJ1t4B9c
6Mkt3qkPqxtlsAwauxs/Dpg7jpTuOGJRg8vjGCsb8A/T0SjuwLFyMrryaCcaHGkFfMg0Y41XzQ+j
dPuoCXtpPVaACcqM/J4G+FCNF5n1EjglumpxgCRa2q0kWzyxTvZAEVwdbx96Y0JugmnzZnoY66Yb
ipcu5POj6jMDmXVaR+f2MQxuWZwf2j3Mg72w9rYaktrNQSmUDyDKj2f9zIXhHuHKgvCCdn67uZvr
M7ibkhu9CgA7JQxwo91L2qJuEFXQsZKcwi/uPbMk46HzF+WNrrUHliZvXx6Pv29X4yR1oy1RO3Gk
OxKDsekOAL3xRe58JbnPSq/nffBnboy6/IjObWf74fafjOc7aNZPb44LGP2hx5v9o+Kdhb7t5Beg
BhyjGZu42pCABJrORlePBuVz9PMvdGTJRMmjm4YK6/XvmaV9E5stu13iNx9pAu6RFidozB/j+0KW
Aj3XcRITprhbWfLBvomYqR1F7uA9vzwjsBtqryflwf3QI1b1E4gt+tR50yHUPD07BbVw8/WFzLUW
UHqzw1ookM5pVUSsmPYkHEnx8lqrseMojspMHATEKZFS+OzOQL/k3dtCB66XbyQcFwmCBi7Rgt3V
bCjwCNxZY4/fQH8HrCmNMxreOivIt4sxZaODWOpcgwbfDug35mK5HzA+nnw6e+66e1wW1PBiFkUV
/iqWmB+Ch2zbpfto8I/y/G2avY9BpVV0yON53NS1dkR8lzKgp6biYREWwCLJcMlJqpy7BSArgLcq
8vWSF3riQgfn5rivMp72m6NRRHxfUzJCwc8YiL3BGzFUWf62ihS1+yFZ82F14GOg+xH1f3GcDqd3
eb0vD6n0Ur3MUzQBIpPXh3WC9vn1x0Opwrqtt32yU1ulYW1kmN9nR8ujxp/QaH1GokcNe0Sgzo1B
14XU9nk6vMJyEmBaJPNzbbQRaFrqvmTCMouhzEX2JTBti5Ic3h57rEu32xMmx7CDgsHvdkdRCg6C
m/ycc7W78bcp5HzScMfeSKFKdTyBTEYhqlTaY1elvCsGnMFa+Fe1QTtJSts/9FRi7RA2ryGiEbvl
UhZD7VURpYAKX0sGpcqVCorZFkZPVZBMC/tbLoOKo1EjtoYseVPi37/GtheiNa7NkTMWj1kElqyY
uxJR1IklHsHvZhGvUgyIPxdPHaqIxaqXLu7RNHd2EEdb4OhORnO9etFn0l007yWFbiOL+HKeesO6
QJmhHygYau+5CpSYwTnZSUfssMYeJgd9+m5kJbAwTy+ATAcds/7A/9Zgv4nNd5a255yVND1iyOsv
K1wbl/3JESIbEdoDlFK7/+g5Am8mu6Qna7dhPB3FSd3xGpA1BekfGPaDCBtu70uALUeMl7ISDeoB
RvL9Z+WQe386e5s6bjBD6iJjOBvQ9sP0BlDLiupycQP5BBHILtOJX01AO6nU8fYgWS1/s3U41AAu
AUCV3FPHOynJZOYcbhq4XLZ/0KR6OZo8A22CrLVkkn7M4Nr7hLvcXpQmsFntE5rozQ/5cChTVoBi
UqvDUi4j4PpgYbnHdhSsWeT3bruMAVC3JZzm8VJoEoZV3xC8ySVmMzDRPkNzILYnk3axBAyqN86y
YIsNm6xerr8RJgiSrbgYh8RrglJ4XGwfJsJ8lBzMrEhMPPmQVhYrxLlTOa2YsCsmiWs9d5lBsR6e
3TgOJw7xFKGL7nDLs1ccQvdx+1Kh7z/AlE3B8CAUHXRbN/rldjdpPgCxcOkC7bO8p59oLps4vlKc
dOtPonkJ41Db32+BUAJVuzu9cjh2DEKeo1k2YWHfkWIbc9Eml0xnQvInBk8tPUDobIQ0kgMerl4X
Kb4SLS3WW9bxDoTil+zn5Uh1YDxSAJoNKCXeb9lnzjExsdURrqBQEr/JtYr7lyRQ3KIon/Q3iSzz
WQDSaqTL+qH2hwn6K74IpGV4aGR8/GGlXdfoZc/zAvAvOOwSpD5SiuQktT0RTnPuX6dueeS68H4Z
RdumQf1ponO4mJvAFGrnIvKy8CVhYSe1BGq0fdUy9ve7AxSSD+NlHFwHPPiWwktNQGpviDkpnFOp
yHKSHRxBUcb88Q8oDjoHHZpLYr08fuKD0JD25BAnkrDquaUu6MhuBq5LBEZxKVwhnuUi2ECJbqpH
qy3xybEOl/XAVTLzcDt2CLxdgs4zD9XZCCt9SAdbqqzGeodjnozhWu8cwilqhu6Jv/KADACG/ojl
kbDns0ASSGeR8HObj0AFMGIhWhtutupx6d8hYmfOEUmO/MT9Yd+8j3WBXxaUiojOxrGROGC4Q9bG
yOO0/bhU10sdJhUmhG9hjbhNAkGRrYVjYy9k74DIQ/Us1Pw5PhdGslkO/6TtFK4PB1Tz/mLrXUKg
FcF26JD9ee8YUZ7v3dzpxH1XvznHzm2jemeQwDdUZRdkaws0wlTzX3S/yK8a0d84PSsi/KliqO7a
3s+QPm9jA1iU4+/TbY0Tqomq4eGdRvL37r3/7aXc6KuBZBSjiymhM0joqKeWyEo3ZgKXdAZWgWS3
EsniRVjEaunKadX1CL3C+HNolLUBkwgCKcDO9MgVX8W4JL6P1D914XK32ubtDsFTiJMUv8/dHvmi
EPHnDsFLcnUhxDEEcORcw2ZS0OmdBfXktVvOV3PmevcB6twezanH+elwdflp6vePtMs5+bC9H7XX
Dv2qWmOuwQZ4FYPSUvE96019WBHON5B1dGcAS8l2wzt3ByPSiyCU5TrxQNnkK7YArhZ1vRoK6qOu
shqogb+HIRHi9x1YExr+KBC+sIQzdNtqdOTB58FFUz/b0o3ukld2RJfT7GjiU7zTGyYd41ShwVMT
WErZ/KK0QMR9mOFyNX0bhdNegBCu5ZW6FjtHqG1Em32cTFqz+PTdkry3lWLnCl49l0/F3doHEqG3
xvmi+loGHPQTdTSdwgpLiOU7fQuDiNrLiuuSKV8J5HWXzs4UrymB/oALUdlySiG2Dx4CpzU176lU
wPr8UNYr+n5FzZZImOlV6t1c9SBs45+FBdP8yCOywD2tOuUwhqsMuEsMprPK3JdHMWykBN/5jDeY
iyQx13eXwiqx1sh/NTUXM24SRgKRP+YJsAcYaI38H1g1WLH/kMx38D+ZRmGH6nfPiJYYAt4kR/8m
JMNPHSTYT/yrazKEAoECbgbt2oMC8hVmL1Vk02TnlUVUNJvwxXFuK60zxSB43EdRw9e4euZ/M0z/
9O28tPOskI8XFWD+m5F7e3MbADbu0MTswvszJbIVy+nq2ZHPG12QFPFHhHqr1NoQmEl9hRop2t+W
AmJP6sdKG4XMLz8UjZUkEEdPNE/bZsEFxLblq0rpSi9hcRQn9F1BGaIAj9xRu8Ge+Enxfu/ZMJym
4RBEdt+JpN/rDZVtT4t4k7aHaEq8ecCIm2B6FCS0eYN81zn7ctq1WzzWiL+bmfyR8BQDyI3L1g78
Bjq+JGGC5zo6Ef6W2+Wjq5svSXAA036iKy52KaODrVMzYvgfi0UOkpRhGS9Rsxt/inuNa38AzuLv
3aDrutMoZoaSjZifjYndk5mKrtkYnK46hG/J0WAriZucQ5MxA6BJqlixNkeUKvPQlzG19FnFY5s5
koMAu7G3mY/6jFWt55ah0jgWLt/0IaY6lK5LG60W9K/x6ddmRhvcrADIn7Em6iH5rWsRsvAigf7L
j84Lfaf1FHyBcposStw8jO6PJklWFjqEFECP6RFNnpUeRG24OwlyNbZVmXADnMPDByKbacgtWTSq
o0X6YN444ceGNyE2cOSTODKKSvYQ3P1y/JlzDwhBbUOn6uYLABfd+nxNPlg80Xv2DQmVU/qGnSKm
zKBXK0m0pe4VWb8mw5km8CwAvbSa0Pp6DAjqgtfvFJEiHJ6V3aZUPAc7Y07HjRwiHcbGyofxeskY
xYkE0GY42c9APZ80RaKwrWEQbjrAG7ddUA1PEfG8/Sp/dRfH7QXQ/qBYgYLvSNOZo44dTcLcQ9/A
S9M4E9gM+mSChChSObDfIK9yjrg3FHcw+X6ZUUkPZXpmCSbOB9ftX4IIvy2W2KrKQaBs6manzAZR
A+6rbAJLRFe5HbCRmYhgHyxPg67/JvJEhIGBOe9LU05sQxnYcvVPuid8+KrlUXcUjDu4ugiZXW/a
KzVGnQqt00TWn6cEPxyXiJXE1CLHY7XPPkNGuXuy594Mx51+KnQ+2/fo7FKsAvH1595CjCzI/oh1
FT5OrdXBMknYE0rmUtM0Dyd74IcDAHXptDwC/rZwVttk6ZWYNUFCqgElY3z30be2lRSv4Gcv1G+i
xg2EgP3QMs1H0vEnhFopF/d/f8C1PIBw5WmL4cZleqnhUH7DipcvlgMVqigxIJD1MMTtthnUnFp5
/3X3PQ/4QFnLnyrFJrmSo8zvE/uKkqPscG+keBEEw81vuX5DcukbVl5dREwZN9sz71F1TQ6bOWHM
3p6WRcE4OqZojC0J0QJDlg/l6hN2LJuDhBnyfh0QuYRLRGbkxmLeblhWpbVE6vBk8qG413reHj9a
BJVGSwvdM8CTf4vc+vv+5rE1s4+ewoEcFCs7dyCqCmdLonDT48lpK9Rwm/TyUTiTXwMBw5u3mrjd
6u07AX4WGqfrXurt8SbozwxvjvywubelOk+wMGMNltJnB8ugNH17a/gfuu8wJ9dfDTwZS3Fwqe+I
mdLriSdVkzA42DrtpUDaB7jivyjl1jucImESxL91Qqob13nZf1OMx2D5RAzwdCLeQlaquRmdDOt7
ghKy9QEFtHsgApQvmO3Mo8gk1Pw0MamZWI4B89Y0NUb0Vpq+ylb1X+ox+M2zBKAxL7hcsZNFgCTy
RKlnr9xFScjjvONyfnUxs7Pl4PPUtX8+lw0bEA83HXQjcrJ6DYREd+R9MvzbrCxcOLScf9yYmASx
WCj1WkJsBYO6XfjSab2UHoBn32EWWIwX7ie0aK8S91UB9+kdcYirjDv7HcxnrOxng8aohOve+/yw
bNHbuuQXYyTgubc/bSEDbTzlTacSPOqPJ7OUYzoWi+XtTXgqBIAm11UaUauz+R/lF7YSuqu9p93d
xulUrQEr2mTPR+UfFA2330Yfr8CjOxIRX+B3K/UGrd01IswlJEF56y/89+I24E42t3XoE9ZwmsQv
s4kh8JB/W7XrWGFh9zVl5NvDC/R9PB+NhWmH+0wUq8Wj0m1aS7QemUqC12Uw59l+Pt6DQmA8A2Lo
xxQDF7d5zBaa76J4/qJ/h/K+tBcDArk6JcEJ6dWvvO2lHm3zotipZunVtmYekzrh+kPyM3AGP5TQ
+DOfJ+sCwhhDm52cXZRnkW3RZMt9kGoRdJ+dWb7PLvJrH+zXf70kZk9Zuy16BvDcy9AFFiUyQM9r
4AD8wO9mfNm0mzcxms725eSJN/umo6T9t690LcIpepcVELnlsGSWr9aqB8aqBv89ntKRU/W08n+b
3tZTNZPvcKuUe/wAIke7yKbXOAk3Kv2QBhYU1kHoLLK0U75H6jZ8yxFyjygB72dD4phainZ7ab29
4GXjd+Nur7cL9VaEsjgwZ/a9VWT2LHQDwu4N/kTCTSgcq4iE1hHEXynh3eGOsdOaZ+SsfsG7YgqI
tfRnYFQyIxjPCkfLUJOHR6xGBXyOabgH0toEFx8KX7+W/kUmdY3Ymti9DUWAnYoe9iWXTtKmhmOc
YLqCPp3tCgTrjogF3rDJ6DfYQBBtALAmBpKiX4L99dosiiTPlVHfPzji/Cb0Los3/CxCIFpH3hqM
WGcfrkpd6Yayqbbs6V2xEFpSZVMQl96sCQcZUQnkNTDzJj6aYFezXxWF6SJZooMCv0QSOmHhwaZH
33huBw4/flppphdJxDVBNNn0XJDti2hKlhs0gqvJJdHpVWiteup4eEftdBqxQXaIhTwiynVIB7LD
U4HzS/pgWM6glYy/hxj8PNpiWZxQ45AdYgNbk1M9yRmB0z83PHe+pq+h5KHjZ8F5RYmYLWUByqZE
XPRfaOPtiYmANj36TBvUfKt3p9aVfnJo5+dZUebx8bKjwLEBTHNPxS7AKD1y7yvZwVVAf+as5QFG
zvASYKHwQ9Y3iX63C2FS4YmmUpiuAA0qfJUc2Ih6ha2Qwguwv56dixHdDZgEO5Iv6/krnGTbKHcO
1KGH0dYQLHj5HLyQPiuZJ8c/DuqpUWbE7lLE2/u8tld7pkslzqOPZB/aDT283+mIgBGhRj0lZr5a
Aq6csfNEGGKnplXiz8Y+SJKYZHTNXLwz+S736nNrOafnLBrHhoDp5hxiMD1hvD5v4ynbQfy83sIw
iLF5Xx9XZPVNMxl+07fU9UCZtRM/EUApkvbfn6TriOZthBdd7QeaS8ZZG8pICeO3voKJXTTaHFRc
rdttxvGHQXnDYCkzzft1W0LEb1liG9wkx+FPksnYh8Jy9kyE09iKmem6qtYijnK1sK5lJFgpG+ls
hfabuzooh+IXxN/06AdtPBUeqx7ltZHvklbt5mEsz8FkMVksQ2U8GXOSE4LoJ/L2mD++eA84tZ3u
k6Oc3O3n2H0gVGJpTFVMRW1t0eBWl7YL9eXuWINR46LZ9ewjbqz9gJmqfm4380G4L9zpnqRvhxYN
3gxukgdumaBqNLwodVR6mklz6Lg6K7lM1CFOcOsDfbQFT88fIQDlth3+t/As23dUdW3+HZv0hGjG
/2/kTCv0bhjuqc4Y0EHqIWDqdlNpVQnTKwRkvjaYEPq+am2O5OeAvJGdl6pz462+wEDXHtLv9RSo
nuzeeG8LI7mvxuafs/oNtrxUJ/KumH8vBbxJToN8i9Onj1ojH6PiLdQGOez5liMBWTBTsvCDyae1
bgFC7FOHPdrFd7KrTwsMIeDu/9Q6QaFHzI/KyrM9jbKafjxoB/vgHAnjaqZEwNAZOJ+e1Vv7Pjah
GZJQRshZKUa8HEJzDK+1uY1QmlgqOuKnNx692MY0xTQuA7MezPtWotx0ZtHBhfkQKs6nyfGYxmw9
j5VheDA5gS7SvcJTwLjmqk9Fg7suAGhSaLCsG+CeKJZTZzgnC/NvrpFk7QxcLjdyFYZgCb0k3SEE
UsBbcE8EbYm+LjYdGn459jBwAKwRmfcy5C5ji1lRzlnRPbvM2LbZZWGc/BuojkavnaL3Ms+ErxVJ
0ryMxMVMRP83F5TvWuPtuTy5nLJY54Ok3bKcDRQDlKH8t/KRUfg5vy5gYCDkg5hWHtx/Kmq8bsBh
1YWYkFfiVikI/qeMkFU5QIEAauNaL5N9QQXp77Ro+hctTnpn51ggovcQdNWXoVeU8VwhM6l61hQe
G10XWoiVeuZ9jVe3TJudE2up/ZmBOgrw7l3w1Ylq1f+WHGpDm1GqdkNMwdWh1RSQWHKNZQNIj/k/
Ah9N4JUW9cyCjGHVXxT99iTNclS+C0XdfgkDW3UYfZeKmryyhRkHAp7kktWRdFqmac0liA3HP/12
S1U+TWsWYiN/E1D74N5hlZuZCmcTV1cF7IGgmL5dEz3kBHztTzHrk+LfZ5Eqlponi0OUL/6nZVqk
t72POB61QEwfHRzwoaCkEX23/83AH3jd0GOUXgAE+9CxAL7ajRP8mllSEiksC0h8TN3WL9tynwcp
ccosO+ht9M6DdbB/12w9kQnABesDo12OGK6TqiwWdoxKn6PHZtT7PkW87a+IhPRsDPD4RGB0dPoH
VlrqToSIIVL7l8Gjawq3jbNdZWmK2dZBMJAKBV029TtimR7KT/fAfsq1RipF7F2mp0EvJskf12UB
LuIUxtWoKYmifjswwXxq9gCjovX9WTWWajY9AYqf/d1jUdS9dRQkjScpStbXjJ7qPVCT5aS8OBdz
Qf+0A8sNGaiuVa25sn9hj880Zco1zk1uTMQmPZkv2KEWf5RlCHDtwW2bGTQIxhjeMmsFkrGWV7Zv
COFBuTNokWvn7mD/4+CB4QMwXrWVuO+5P2TqYgxgK9PP1EtJU7H5BhuF/JKg6mHjX3ttCDELOzAA
x+m93jMKwhjkHEtUlqgs/CSmAnFMGd3mQbDHKb812lS79tXig1Rn3pq2YOJdUC1onFY5YFlkx+OR
Y7auxt5x5ci4h4wyziQ2+qsf3G2iKoF0MdWxqYQRKGy2D66y4QQp4E5R6yBFtlSUa85rq6q7svqG
TWbuLfAuCU/ZjQ+fTZuPpzKsKjnkK5g33KeYa1g8sbFW7Dc3LlUKaEe6lIPO2jQtTiEYGYeungVA
1HepKrDjo5O1y8vFw/3l0kDslriAskMXodZuxMpZLKrPyDQCtNpmGFz9TjRreKpWUYFMqWEvDLdo
Z1BYsI3yrEsBHc37Bf84QLrvj7mfAMhTMkfYAGrB6X1S3Q7g74sbk3k197+u5EnsJ0XFjvJDEG9V
BAkFS8lBBij9WnaZ4ssRImjckjEBEil5d3Y6PyQZn/qRViHi4VBIPc2gzuq4KtHd4WahxusZBs/N
REJC5Nb01LnulyFPDPx9ER/HrBVv5RFLFmsPD4nuo4oTdFZP77B6lUOK12geK74zuAsPwRixHv5N
YLG8xQuPY3fK25w6fs6FxpeXhESC0SuAGlKWzTsvAMymVKY69Z3RODWGyQT39FcVCB8P4jr12twP
TAPH+R0OuQONzFhIMLD1EOuqJz5mSF2xHHLeEkOohpAPo9mtUE6+XJXNU1dtWYEnXtgZLpXrIS8Y
qqkqVP7QsJzyS6qbibtuRvSgbbVQ6otLUdwR1LaDvUvMQpQoyf//FZ+lGiR7kMhxhIlbSj7ZQyJT
sZoJZ6q33iznCpMIhH6V+OpwGGo79BGYgxpMRP9ZTrHjbX0yfbszWtHeWXyz/gzXHq0oCTTc9w8R
8qvgXhmJa+xSh4cjirK4qY12c6lxVdqkanZ0YYLvjSNWK1N0wupOp5kk444jH4hSNcYgSPiaHzj7
AR5rUyKGhjjpppI1Jl4pgblJoqJ1k1SI5JCx808ym2X1lWDa1jNt8PCmLxN++/OZ1PbELx33GK0j
8l4fgCmysb0WvfmRa+uNAr0Cp4tUxeLK2gsPsGjJidcYY/C4Tj8vvS2HLfFXTlbmN8UWuX12SI8v
GJiacIa58VJyPyjhfvZLl17zr8bp+AlKAKiZcC10VsohZiIM9575FJniCdE+Gs0ChxS08WRQOegK
S/oD3qAWaHt/eJRe07ilmbajG1955o+Nwb8xVlBVgzvjUQMD/6Bx2g7IaFbJAVYSZosar0xk/77v
MHIyTcbPEXkLlGXp/dnJTFLtmtq066BjsxQxCW9iiUPHuMNdxfOvdXnA8EMZxBq9Tsnw2c1Dpgto
VunMDZaant83GjuC7kgWxVGwih56V//8rcseYSH3Imk38MlFOJ/KNvqfNfjY16X8Z/0HwDBtfnox
B/HJSyWOr/PHZakZJ6h4Cbn+v2FBZy9XJIqxS4JB7wDpLyOn7Ue9Cw+trpnK8mJjywMaYNxxPU5k
QOQahmc5kfUNlPC3/khR+S+jTm6GG0ki2RB/+2PIgEtEoWKuHfSTUdS0daysooRlrgZtpEyPTNXu
xGM78Z113hcEaeSo4c1NtoVKxp1ite67Qg2bhN26Ph/NWWmKnB9f3kBJ5TKSxy6Ni7aBF83RFMYx
iQw/a7Qf82wyOWkpfKMVjtBVdMh1g8t2BTGmpXAAK+QpRSm43TBiJzVQmlJnYun5CI8yyqb7VtN0
Bj41qpsVaq6jwgYYZsnHl3BxgnCyjRhRQBvPBDJYnTFAU222BBwrQJv+CtecH80wnlrahM1hu6YO
aT4F7+j+EZLs0y0MSecKKnfkx+d/Ns+DaXATMk52hrlvvcoNVT2Dtm7rRX74A7cdhKX1B/tLV/fB
Y/cO8e+GRnWJGz2GtgBhniLiM6LQ+yHU/YmSJrvvPJNqNmHLXoX7eyhl/b1TsZSr2uW4qTq1sg4c
hovbO7hatYsaVNx2R98z92DvnstHd0uRtwGLuS/+5IEdhm9AWcG2EfNZsof/mWEOWTFe8FfVc7Md
aMkhbExbhC+oJO1eBq1vkFHKUBJxWrvNvNG/Q9LxAqDZg5E96GEMdRn7s6c7LgzLuWG+dHjYmJQk
uGzZ10yRAUNxIa9hBe1zVUwpAqiwf9YBHXQN1zYO0+q9bHs0Xmay4vSfu5Ji6f45F3f/WSIjPV4N
suh/cDemn2pKPyp9Pjw2NRGE1SriEXiNWrGKsVckRHSBBUPEz5n+7/dHQqHeNL3lNxwf4D7xnw1R
BhAi609x0F5DPC2cWwlJ5TAyTSD+1quQf1OFVyBaEM3x1OaAabnDOwGxGj7h1+oL3wtJWEgJozzo
/iwE9BqxKZloN80jSCZyuo1WriW84EsTTsoXhomo4ZG4aZVLLn+lXZqEeLhqSRDG95Y99i5sc1cF
u0OOl0kgOHoXwIKdS9/ufHir/mQ0tcnKmsdRWG+REq3+5QOvbj0csNfLfiYdc/scEZ56XE/qlbcb
BA+Ew7jwbHRIjB2Nh+MBmJb385MGKWw67EGrXtZrrdEboj28jOuOlo3Ku6g1VrTaXEs8QGz5EYyc
17XP3Wl0vOMz8L63fWVk4nrOWypSD2/1kzwkjWr+fZY0rU58tPv0JBytagcC57UP8jyNrCHYmvOg
eyJQAsxBNbe4rmy7k24IKGp3jtaqSUe6qCpvPAEUjNja/et3qnizy0h32ANmsmCs7FNFpxGnfarC
SjEMGEWtWRo2npX+BMsPKMqm3v8vjmhpj5LeamRyaH2cg0xi+NTfom3vb8ZaTOc0RjZZtBHznt0L
mAlpyArWBBjc80oopeL+n93yaP0eveOJGjn1PK0Ty2ao2THFxK0B0Se+IWAzY4XMj9CRpn8zYK8T
aoGyM3jJzJBynHzznspWRft5ZyZkv5dxkVUNsIfGqPI0qCQ384/2RsO0Cp9Nv7c95uVjyw3FQ+5i
4uxHmRfxGIhJxH7+affSRWFAoOII83tTiwFzRkQTYoWsB/11Sk99wwXpBVI8rp9aAQSshqjRjHak
8CWfl4e5gi/BF1V0+j7lHmhDaMb77Bi3MKP6zHg24SXMI3NKTkbIMRLBU6NvsO9RyslY93aePh+A
DPhCjI+rLEgJlNItsDbCKN2cPyTCHuzrJUvwXlhF/AsS7IvcLDx/+UXfhTnB4ZsVT43jbBRkyVPe
4lpb4esr8nzY2wuOQJnKxomJ6s4PnmXUoUjrcxo9k9N/2OhjjFKAKJmNs8UVjYponp1Pov1s7zWB
7k/YzcU6OfPY9isAnBGtPjit2MECECm4F1I6wQ4C1w3BKJGs8MIWcHf/RWI+Ga+dqie3q/7t95D1
r+iRj0pXFGbJh/OpnZRNMWWA7w1cav6a7Moz5LOqS6yxcG19s86EIsfjlXW/h1PMHBS35ZHB37/J
jLnOgsbYKjYp/68zOAFHEwJXBJE0BLvi3iwEIZ4TOAAfdgZxL/ZDIJIKK219JpHJrcpmoflA/fpp
d/00VBBNQcJixdGehRr16A6t1TUwxnsgOPOeU0xdl7sjo0olMgR15LCtk4dfuGUvLxty0eFq2tCY
uVU036OAfPOWqcI77u2ujsY2fUlQ+A0yIoQdbYnUcex+opPa0+EWvAr5V4KFSOF5tYnQiFr6N7eB
BEzi1SWxKW3J37iMDjeRqekKiaXEbtEdjIV30pEULoYC/k4uXo/hb+OWgNDd4dIoDJpr6tp5poyA
mqmwEePNMpgwttPqN4fEmtjWufkmYZeilOtRxD6f9SjK7feJX3WX8tTdqKjm8ReSCc/fAHT05vp0
nNnaKP03MN2yVu1h1fdLoS+ooYVw+gz5LndAPcYkGSx/QQKNsEXJcBnW707Ly6jXO6095bm0XQxv
eydnk8TdGjCiKFtgkRQQRycNoA0Yg9JX7FkDXL004d7gvbK+M2yQuk040bWfTGBulNWiczynMQoU
2FppmHG9xsFnSSjPTkHoL9eGrTNk7ct1sTC9csgEl77aMkKkoy1ggW2vIgr7w6HNkW9iHHZNDagR
o/MXC+3Er4S5it6AabGM8fHFCE7G2DRazxNQU1/VryL8GCCmuyWok+qletwb+0I9K316lRzXWrJR
gZHfnPz8WOFehVKPuMJ+QH8rUwRSasYbi9jEcIFXzH9lp8kw+nqtIDt0ulajRUbq0gR9FqrVvlYF
jO3PRL+lhoOWwPHNGn8NOOxCAn8/lbcIcETqos3F2/zKoKu6gxRM/s8LHgs9lPsjHFw9f+6TJldM
z5gRrEkhRJ8kc11dbj+IdQjhXtLeZikkmxcWEngpa4UDpx/WcESPoB7YHmxSCaIQvv8YLI3Pm1U9
P0fIWxTtAwnyfpCpvSoy3ARh535OcEEcaLHwoHPek13H8dqrprLgWWUbkgAtkWqQ2J3lPGXgm+k8
eCeTo8G1IHOT9Xf6lbVwmJy2AcyVqZr13kXGzcZ3gO6EnLpzXdxWM3+oSankTx/O9YDIMCLjCISR
e806Fi+RysZ6c5TH9LHDda4348HROj1tEU1ik+HelsxzYq2G/J2e/zR3S//hrcsynSEzyFztQ5wT
K3RmNLDdJ0yIziYpCDLNqALfXoDzkLEdQStKY/W+2S918/9odOVEsoe7vC23MIeNTeZ8tIjRDdcM
bERN/xMnJ3Ull+80qm+XRn5Gxxn/7n9eelNNIQqTPEgGxf5J5/yLtfz2lzQmX+Ke+Go3Fh9SZWb/
Bqqt2etNrsV/Cma/7g6g5aU2BnFAXbzsfUkPY9YU0ZL4Majg9oapOS7JMbasjxcUGT4wvorr26aQ
Jkni4vm8+nuhzIcz51jJGVDvWdulvQ0lUutoApoKIryMRFoe6grcBd8dmuCtrGHKz0buTAVS8geW
3M8Dmx9uOkOpByhgRkuDsqLaYHk3yOpowe2fOeylQv7CrqxGqkVP8NCuZPhpLLNwX3FyzpE3lFB9
efoYea9DpihxIzM8FVx+3tSJnxXB0/zn2szPhj0QnqftD3VF6A5zR/Uqrp4irSAHgO1Z90gfOmyX
KY8FDmLRh91eKBasAlxAkWg7g7leZti7mCWMqd35EkLitphcJsTdBmSAsRa+a7VGsUo06Wy0DkvY
sfIYlZm22hxD5X2jKQ6qACZucDbY9PCYe8Olil9BLmQHxy7qP36Ctfq6tQGLDanzunQoZ17yZ2vg
Oc0Fij7MiRguKAAD8HPduoJdzfwPj4vxOxCAAqRlVUsyMkPnBwp4sQYQU4th5zUfXqofMgKfYrPw
j1GvyFufTWdsha4ry3aoUn5bmT90uVey0GCOutawPiBzIP1kKnZ8jqPUVriTZ5ILTwL0MKqJ+IFk
eqvbx+/X1KtcWneTWaYaGyOTr+IR6gi7jeJDZpX5xiFgn/6K/A5iqHbPZ/UGj2vhX/Ca3opicee1
UlaRb0GCDOZWllL80qDDkJEnBb3ZMMQN/q+iYDq49W3tKS2E34lxrS71ILPk1SqeNZ6r0D3BnYMS
gMQYEhU/ibwk5iLNM5C4PIKPHi92QrjR8AD3fCDvIeetFHNL8fTUvvDxl1dQAli/TBUA3wJDE2JV
GH10fDCVo6EABiWng5ulIYK5+mUkJolvs1rxinJZTXvFmCvjXa6zQ8SqK1QwCr8bgjFONu190t8q
D5KuVE2urK7380UPr0mC+vyg3hDhyE4iSQmDfjzN+qTmsZGvGG/84wJqY/QpCG/I7A7WNNrmAQtq
oec7m8zTJL70MOcSe6UDc1iu5n+TSmuESwNDwzpE2qW96Afr4KeFpJXaWvk/ITxI0slc92/SrqBs
5gy+Z0wJCATxV4ooYC/ak/1lY17WRcvWfEtnZzU92vhOJ+uASHko0sHNq6Blh2mTiynTiddO4SAc
s79W6NPU9DPMev7U7u+6Iasea50WM+ULdPCP/dC5Y3bbnLZoen46qyRVQHj4pBqzxJN0vn5qq3H7
ziUKJRgJ1HiSN/9e17t6zEkeGpUUQbzCRynKhFXdOE1eXjAcvHREgrtLQfAO5dhqxcHa2IV7hFJr
o7N2M+3uwOEKSbu4PWYvIpxBPcYXUKgou+8HGdyDIPrcjWesCLiscO3r7FQx5NUE/u/Avhpwy9pA
0abAKcZny5ssvk2iKe7xdCaJUrXlRlMWTRyyv/jqXRpnmt8fN+4Gf6Gz0TKUWvvqYfvRLPjD4Nk8
xDlRCpTHvXHmZ/rPG5iOsNOGj/3+SVNsrRglQlP4NqFSRUV85poXUHZvbXp/qTYdKXPkyAcenky8
tuOlOQ9TfTMtCnsgMHZxT4Z/VlPFuVJFxFMtT/klOxdqWO0DlGtG9BKDyvmkb5PIT/DQd5Gz03UW
WH1R7TvW4q6ca/tlZV3TzAUVe8Xi1Iv2YinvSCitaHHqiWWcX8FJ7lWuoorPdY4XSuzt5e80olq2
T4mmZsJwOXOtY78U8n0r0xncqNFr5JlJALw1+VZH/eMJqJS3eE0qJuYHFsX/Zpf+QKJJj8vKBveQ
1DXhod0s7NJ4zTs37z1aON4LT01CE67ggs+ljd0gKiUPkqXxubbJXPpvbfQKPEyeLeW/KKAe7Gc3
wMpNZS/Gn+jEgdHxJMa1wCrZW89bC+iR1DI7cDUNSbdLqavp4dqwLLRnPZOh5o7NSDhsIBY2HP5p
cruHWsVTljmcACfH1886nJH19Wb6BZjedeA+vpQL/JZ+luQBLeWBgMqzE7iSRn+kk0wL6zmBpUjP
xbe5BEQ2VKMfK3ASLkU1wTh6lJORu3BLnXyEks7gXEjPaNXl3QbZPxhluljWOYfnJ7er2+sofk0y
M0OfYHqGfiLHWFiSn8fV3JauHSsqwNFIjWYNgIvbNG5aAWSZnuJA7k99MYzSs9lWLt33kX3wC3xk
dL8MpEuRRvwZMd76Qk7DYZqSAdqPbJYgzFgxj6eCzH8gImM5Hkj84y+CMK+tYXccARYVPdWfuuyF
w+5S5hkdqYNLg7FJpvLtFNKn/ZaynEpK7XcbY7V/+hTXOv0tx6Pl0zddgVvQrYO3Pku6r8rsCDCv
rcIG3BCy9632PHuBRD7ndMwuGErUjbC6HpnGhS20VhgKZHwxjnErAjcVskFOIe0UGecZgOtTv6U3
B4wGFj1TiVl3pFhyt6HN1KMCS5ZiVUK2WHavib5ik31HYEvCPUpxmtR0qr9rx92bV1dn8NRecBTN
Sbg1I5QgKDyX0GNn/qvR31LUMgrnBr1C1tfhrdKrmsDWU6sYlv9FP8H3p1oc0QxtT2ly9FHToHlx
BWn1+U7RcQLYaTc9evsPxJ1jVu9gI7g5Khw2Tn3TA/z3MXuvqJa99RKfV0/vuOJzDcT+DmlcC0zJ
xNoRR2Z9UVmAN3dt6QZqHNrhEVfJswHfJ54E9jJgDO+QYyGFqu68KoE/D+tsKumPHpSZwN1R8WMH
cEG5KueRr+E/bkqwgCjkeO3QVRPGxpar/o+BELxfOBMx8U90KpssjPtag5Wc+SYfvWPzWUWdqYj2
z25zU678liTPYDK8jVOT4cjZj8I7H3IC+4aoEokY2n2n4VRvERRlOcPPjakdc/yEZGVHV3YPpV9n
wcGyU24lIwLWiD8CxxnA918oKSr3YO1MvRdaaCwZy62vYL745bTaeMctJ0erlzIegBzk1OaUl3Uk
0kaADIuNCUGOL/iTrCqM5X1ImWKQxQmqziC8aR7YJTP6chcmYWHQJdRVxseAnFoCA9OJ19j/nw/f
eEBkX90+o21BgO5doEeWGMC49ivnAmH75bV88u4fuh38ipnCpt01NBpoOvr6SfMbgO3piN45lgjp
eT96b7eqXsu9GrjzZ5aYSvOmEAWipiMPW/aCGPoaklL1XoFJgcE5653eR+hY3fTt7VZejet/N7ZW
CgmVXUh8BM63sXkYYRcQK5PRxHsuHe2yBtdlPCOxuIrD7EUDZUB3g5aNd72zygYIm6VoLKUVEMpD
LwVd0hoOpJVaKZs2Zey9391bJ+/YmspS/a8MluVbE7Y4iyVnu036kTZaftAIAua4l1GD+mHb2pQ3
EaBZquIxHa5VM4YOpaCpFOYGvIRJaNuT3koAbMJfh+tb437Fq838eEi66TiKgVjj9dFXXu17uVrm
FltFS7N9ltTj9jm0y9L0wAfPmlMePbGL7L3x6k948uT+cThyrA7C4IWDzzDlM/z0ZzHkds21RSbG
1QHeMAvGXGoVd9mc0NZmCJ1wN+hwXKE3kYASD/vdaM90K5rx09eyYRSCUYhutInpvQUYorAi/fov
5r6EexTu0V6vULFVrt32iSE7dZUns/ptPtqrQfxwkV/CJcRznt7ebmsG26pMPc/6nu90dH6TGB2t
wq6vzhKtXbIzKuCRcJCYQcr45z0VRA2AxU8+t5nZPgW8DM2sSbdPlgoEBCGVnNVaR4n3mEGf4ONK
zfkvq2QB/1ou1OXULW6cwVthuRBPQhQYmTr75U81jEEsxRpaSmDjFJBTI6dxVkfUJc/Clsr6UwO7
O8VFGY8yjsMcZ8lVpe+7NpOiBGqI/z51BaXx2H0x1y8NrmvAQoWqpk1xOmJQc+OP7xWilNn5ISTF
QmZtKVbZolDYVnhBpMp4BikVHbAhsUfPF+sTywaW1oelpOrISXVufbFvhUNgz78RDfV+UqWMe/d2
pRsno3bpagotOpb1oWITSy5oO/iVbAaWjC0TOnHMfBP2gnT2gUu7RqBmOtlDYOu13ahNPq1zQUyp
RaeWo4DQC6JgH7TC05141mX4IBHWib7Cu8w8G4aN6EDx48y80QzBoq5t/iFLm6iyESe1iovAElqf
FiBStkoNWenagoz5WAresl3Z6BpP00KPa35MzbBNhokymu5fabxGfk8cK9Vsh1zh9nxGxnkwr8I/
zakDj9t0DlGJ+6gMX+uuVAFee+CCBUCo/8DVolfIQkHfFGbnogO69tewOk3etaNSD5NScqYXIRdS
BRxAQMDqUnludjTCZZYm4vdLx5CDunlWvpB1HSqNC7ZWkHlVyKgvaa+ImXV2V7jP3uwvBQvr7aXF
WsBN+9lHl6zlPSZCA4hPzHvv71VgLOmWHSmzRzGi77+gPqmwVOJtN4pmUCrECrNHIBSFshTPRs4c
44M/6Pbx8FkNCiebfU8f1v0pC7YWciqbUCtL50+vSfa+TxEZrKJ/agGJB1uYoYfVFUX3a7Ur3YNU
cOZx7SNi9JAlk/xghq3doxBqbFA0OhVpcHcaAIfHF+BJujjOQIl+9q/fFhbhAsc0ZSH5k81R/SpI
xjcxb7BFdNW7sIqSRqKClkVyIckHhfhhpKXcFS2deMDqQimG7JOHLykJckMRxtcKW4sSOeoop9uo
xV0FKCYwI5+RFfquLuD76Mhew3E8C4B1Bu43uGRvIN4r28hqMW1OFml8/+hRUD8ocXwburVRU9/k
u1sUktREevEAXhzN4kQbbQzBGd97So8dKrU2eNJa23iycZKy/+4iE+nYngtr0Su3EHISmq7cEXUF
ngkH96PnAXartc+M1obU6saA1cETpbPxddaECxY2Wv91zJ114RlOq6oCOY+ICRCL9lpYj89rDQHn
AgWrINItXqtQ7tFBz07+Lfrf5bxKp4pIYhVlMJX4139iIEaLZ7d90Za8PrmtyHcM9KCyM63sicVX
V9AZvMfHrpJMutOC/kkt0k+Qf7GH9se5BExLLpOFnQlDccs0P7vy0p8zNimQmFyk2jKSaG0KZmO0
XXGVYHvKXNU8uaR47el2uD59ZNwHq+YU96Rt8t3QvibaujDBinymVfjzSTj79spqmFayToq38yTi
AmsOtb9pTplN678cnO246qiFF70PMOw8bN3lx/tL9TpWlERLYXzWzwhQVSVg+51vHTEb/ROQ3MyV
eIiLuWV4pFEBhnrpkS08dgiFmYtCbkUFVCHjxEs6Il0ruJhPsWzKVgBqvwGPSAUfM8KIW1wuGbAO
a9Bpt69J4UHIvV/heYcyFAxEBS4cphVlujPkkyoAaO8Y6fRrx18n5SART6TzCOMYc3mUK4ryl1h4
BfzqZIWAZgR5sFulieBlbEFAqdSHUh24E6aYifAZmEv2f5fvyLPzs7toM9WHXRsP/DQMwhTb14PR
GSB3dY127LcC9anaGKOMx9/zy0vsZ0T5fVECj/5SAlyW060QuzhI4wiYo5FOhkJdykK1WBYXjNOH
y9ln+Se0xaheUN4+n7/2N8UzNxxai/rpa7Clw2kDOr6HE2ovqbtD3ff+R74OzEJcza5h5qsQw6XT
LKh1M8gvac//AKx+XZknO9qePnJHsXRveRSbj+7zrG48JGKgc6+d7SwuY0x3dNRDLOeGQqGq0GXn
LxZLatL/moRotvc0hpVn1uY3OvJ5tXZmEm56tu44rL8hs9Ic5Uw/dPO0b0oy/pbZXe1v9T4BW4Kc
48X9XeScnc1gviYCX5NoAnvYgvAmre1+wJwB5KlPg9g1nwCarjrrHfCzrCZWpas/SG/als9GeNVF
r5qy5fq7DwuXxTAIdG2MbBQGNlnbk82ke2uM9qI/aIlYrDk82PemvCViPDlV/3/QjrskSB7zsQ4G
N1kC44w8I3O+EvJvZu82Wde6fP51NpJ8jvn5HhfEqLep7muawygni5s7TLgMmLegxMt7XUYwkt3N
9G9Uq+O2yUadUBnQEsKdbzHr/n0xQmCpLzq9jli+uriRsGh6cWqYvgCIhkd5VN7RnrND4IYw9uIT
h+RtL7SrnU4tnKvhcznd+R8R5krkoi9Z9PExdN7H6zp4oPbbYiRglCnIIiFHdDNGZzNWJi8325/S
ekvbyyV3rJBrE8tLCBmPh3t3zGYJJTIHZf4Yvvdoe3w3T9dddDM3eo6Z6ZkNtfpcS6ZnxDPNyiRO
qkkqv8UsG8c+5GhzWr/7sjfrakWus6lAh3CAxQICB3AiWX9Eoy6fvRimNDTzshOI+nEkBw15U7nH
Z6+Af1Kgk/1sYMRGkXwS1KDDAulxmEQSL8MakWR7OV9XRf+YEWFdBfy3CGOC4KdSyQCxEQJ5VIsd
H7OYOfMRNwJQbmpCvKfRoLuFXDsSDR5ZJadQnUdylbUMvcn2udMXUHnKIPcXGNnZK32McfnJ9ljJ
5vPCPKGjP4hQ0YLr4lmGQZAmY9OP0PNEcWS6JnfIzGYQBsPW3MRAd/p893A9saCMHkJ5QVtkm6tO
DldkuXZOyFFpTjTHydI2iR/9jqy/LR+wnK7tfGy25xN4YRgGNj8ORmkWX4Vl6WFh9AY2NOjG2eSa
xz+Ft1n8EoivabybOdzZ9AHhCmcT201ClOf1Xv+Drqkyrs+NBL3IQ4vZOAJfT6kPpvWZPaKnLE1t
0lP9DlCci+SrfhMRzS4wdVOG4Xd/7AzcCp/Z01RcqmHaDkV8tc2JvnaKH0eqwulIo3pUk5L6kWyR
bJqTiOH5r5x5W4jArFQ90EfEV2uqqOvNgQ3h9HDv9Bo58epQQhRMdeokUIGjsqD3unXwdqbTztLb
tH1g8BZMi4wSmPkyNzGOPbP772pgiG6ub9CMcmrBfkZBnNnHcHO+Q+EgsOSahlIBbZHxSXEg0ALc
hLeRICc8xp0LrEXTuAWyiofIH9kUVMkCNldif/F+ZaUlp2eBlDo2Ve0xS6DZtszx8yo2hNfEA9sj
/d3FykrSDXM7N3bf4fTFdUjzLKSbdOS01T6PyAyz3khXU3u0oi+vHe4ir06j5etR0+azGXNrLQdf
DAn6UMbstm4aT6Ofyv1iH2rKpCNBhwDlGGc/ZN2YPh8OAbjl2tpGFI8gtacKR2v8uXyJhnnHZqDu
PPCYtwuE8ig5K5zBGG0Fbw2wjk/B0wfUz0JOGietidGiGHGDmntMc7wQ0RK1Qfex4a7Q7vIlUPeF
RVRMQ3IC5e4yBAnh518xg/lU+ty9hP+rMZBC/94HTdWpaIQR4NoKu52sA/8hjRDn/Jq0DznPyLyO
F/AxRloI3gMlzYN5bg0P+A/21aofrxDpys8ljvJrMIrII/ZvO1K7EOjAyGsb21/FySVENAxj8cfO
LWz8CTzn6pN7x+eH56bBYfKz/bc4BZH3V36hSOCv693c8y9Da0UKpwC1GW+PYbyzV4nh+YSyU8TS
Db9AqgVmOZ6FSVLuJZgYRPUjSdz71PG3XsT3cjrza6wqPEQIK4l1tdtqh97PlpGbSQJaAeu9d4yZ
OFbhMELgIG2GBQ+Q+h4yCyf9Wku/lEffSDp6jMCJFgMvTNEiuxxxcRf1o6VPR1wqmeBN0q1VJYtc
EVsIkQXpcrRIrDtjMgg9Dg6YpkS98wjP/eunCRpM4HjOiOPR2spFJxcS0RHqiSUY38DgXV6ffnf9
Lw6d77gZeXy0a50LaGI1qsnaxeUV+4+vkTEIvHOmZtp7Cv8mMTybjM75l28WZBPm/nwUnQvbrguy
fjIpyD2NEBzKuv7ZMCw0Vufv3QeRjKImtsNCzHliBrsYKDfaPfuf0h9Zu1sc5Ihp7OU3Acoadkpq
BxFbXMx+LGab1vE1aIM87MixyNd4fZlN2n/9pqFNavGo+jyCTrtkUL5/stDWpXb2hy4JmPD+ALD5
OQZjoqRtE8MsLzHhkLUbFJGbqEkEGzTyops2bgF/XpZBRq8y272vgYzwp+zQlPAK3i+bXxxZrto7
buDdhQLbF1SPYAneSLHDV9Vft652atEGfTaCI/WXB2UtNk9Sks8rYY/mi53aCQOnWk8LdkzkW2rv
8YJhxnJ5m45Y0ipg5UCpB2d/oXtxpSsZcxXCLsJJuVMj+vvAX8s3B9+28xgWaylepV8pE6k3+d6/
V9mXXGXTdydI/VKcCs3x2Ya89cJZ/sZYFB1WYn0QZeiLFv9d4tunFSxEnaezSW3sx85EVsqWrgbn
TeGqwJF99STy/UAsqMs3HhrgLQXU2O0F/UAJ3saIDjdeWAgIV1ffaQgkZt0dcOqeoY1Hl/89wvnd
oN/Ds1goBSjzqShotNuw9d0hUPDiz+wfI3QFF4IEOBMkBmyf+amBW1PS4thzPGG6WmfIUGFaY4mC
kahwPA4SW916Uk8sPiWq+0EJ5BCF0WFfZSONReDOyNQ73//hUjGav77BcM33FaUmi74IWFQvF+Rt
h3AtxHWR1v9tNb+YwsW+X+u7AQpabcFO/oRUxQcnf+VZJTK/Ets5t6W1jCd2srQf7o0+3NaxAxM0
VswAXNnHuw7VzxMVSlebX8qZDFX8DXTWo+zd1zCCZ1tHat1f7reHNl7jc1yMxG+XdQjJAZMQmJnq
65mYqHVUcQ62EAm9QxnTQAqxjDp448505ioZrcLQiD90Ivx9C5KkzExMRO7L079mX35mE0gMhtC3
OpyuyDwGkjX8vNZJ/w0fD4YLamEvo8yyV3rsuVbl1zjvy7evYFCL+xApZDwabfqgGDBytdxER/Ws
iJGCceY8RdtX9yuedZm+HpqDu001laVBhh8FDGgY3d+nAZQiqnLRa1HwwedFcZHjcfAGOZyX4LUx
oflWmdTH00eJ+4JNY94qVodL6NE5qKOzh9pkW/8c6M4XEPL41krm09NUuDRBdQVj4FXDFF8/m/Cl
PJtPoHpNojRjkveO1imavrF4pkwuAkmuFFf6RuNc7Ki5l5iJrWrcgOX8ISJ9AVsjc1ytsfC7fUQV
Ld/+k+JWW08hwkJmtOEkSmcD9/BZxRHZCJSeIVfiRH+kn0WhgQX10pPM3Bb7bSO5lXiciVOSuVCy
areh5kv1t0P12PKakm1EvOQByFkNM/zJs8YYCdl8JzLP4GNpc2unK3YLb3amU+ubR5bhW9Ci5YDu
dH1CP5bXF6RA7eEnfZzdeHI1N8O3I8/H+NtGHNMTZrsxObfnXDses4zlQigne5iqKp0McsdvdMVW
/+olMVab48rCA71eNXSBWwoYfTHLnTjFTDnaO2XkqjjOhvjqQNEbQKoHEEIdcrsh3Luwgnc+uzfg
WAAPSVeoB8gdpYRGV3csvUYq+vMp3IPqcDKi3gPt7cvb3vF4cTr2Ui7nQyojtTgcDGFEoeT5f/kb
ttoA2t3aszUvEz42fyEyBucSooqoISO9B/3C4aSUYUVBcyRRT0Ds0bB5L3bKYsrdjaADQzxRNyQM
VF/FyPR656W07TdnSiwFY7XsiManLE0M+KqptWGIfYbJDT5YPZ1/AoW2pFpc6pJFRjEI959xqjPo
/m8D7aRHCzJMsKBe9OOoxVTSgqsBvdDqrBDs5JgS5MmO3UKhyIHbwHbISCngmFc/GUUL+UClqeRV
doknGfGnfKeUf/7Hxf5nxU+f8r7NXzlZ0IsKb+D3B8TIMZ95pQYMeiTOo/S7ltMGii8XXuAzuNvk
wGH4KAUCtrUhw2+F3ldA2U5cAjso+cbmf0gY4KCEDF3T/IXjHPuJERn1rp6ePxOAxAFQGTxR3FaE
+2gR/eec5b4FdiU1nBHhdZuOqIIpzBYcwYIjL4eN9Ntff84UBCpRvjB6GIWZq/LeUG40pG/zZro/
RpJZH0pF3G5JTMWBo0157/RBP8iTUo+pT0qvun0E3cd3N618xoGL37yhe3JrXMlzfMIdWxpf9By1
s2JJB7URR8IR3Vj70nAJRPAApUFefF483CPV8IpYzMvUtIn7wavpttBsCHrMsa5EQnRxJe8TGdEG
IRr2w2RR6HchsafXsf2FOzv72JlbO/5p57GNJp38PAAt8QfEg4NZPQfFbCtRjNGwPHGqxQ0cYCEa
yqH9rHm1DCID7L5+W06jvXhZ2CeBEv8oGyJmOGODCs00QWerAxPan6r9x7A0NSbUOB7CjMSKs5Qs
wvO8NWRnJ/0Q94O9ySIpYepqFLZ5yXoSmVlRcV+dBs28mL2YQN5DNnLMR8mKISbEDJc1dexlNRIw
ZFD8gRieSnP5Xih0ZtMeK4lLWYTJUWf7qR/ggd5w5xVIzuXf1OR8Lya45qMPF+SSAGepfz27XPWs
q+485LZONawkhcu2vWgh8+RpAN359W61SCx1KiOacKH71O1Dm7CAqlkANvfogIofbiWava0j9b8i
exCwKQD8el/F2BFwNRLBKZyPPeCooAkWGU3KQsRqEmzFhmxjphaRWfK6ps8D6yTYACGZrfS3hkP5
SMQ+JoUks/SKY6OMYVCYOtr7CJOQKIt8XJO8tSU5PenZgzSHV8gT19BoUIxS6ChMDl1deT7/lPNs
fFc5D7g7XfAus68840X9FZjWxblaOUIWk10PP/bDLsUUZwo1XuU8f8YVqyTRTGSoYI2ZIAe/XDb9
4MnHRx3PZIElFmDlPiXhohJPodRiTUQUK8Gr0QcqPf+VGG0ADTjNKbWBzIjV2YS5MTN5t/URmTJl
Oqnca+7abILCCIsRqsrIE9hFE1aLw3eo9CNeNIFhj8uDBEGVAr8cvpO0yl8onhRu94wmhf0iBhxw
ossubYCDX0M/bKP9pGxDY6kL2uDrXXOGXlCuBZafHKjssXl5VLkALj4XH3fxl5pAXoLuwx2ZK71L
Ir7NOPmSWSI3AeZfxCBavB42Q3egQ5Tiz+kc3QBkJGEfb2asXU3g41KflOu50fm9XBaarmXLXjmQ
Znv+PYdQWsoSoC94V8iz86AberRqd6WVhWMFxFwmWskM9VitWVsuDmoR+ndOWzMd48boES6LpOsu
ijKk4h3qGRjWl2sCbYoY0otCHP2sQ+BgDKyL72CzmfcewbRWMdBGFN/c6a/MannuIOSPi9UjJzgf
ma/hOeU/B5K54HqZf6gmjAw8eAAhH8HLKRekxC10xcuoRKoxTJX9ystdn17i1BbOUIcF+r87S6JA
vaN6a5YZHSkPikryJcloA1cEyqCTP91ZJMJXtlKOtwd/ALgvyf2Pc/I4g9Azp98nuWLWZBDgutrB
JRLPBqnGj4AMPKJoKLDBFLgzF7v9NpslhjIBU7KPjT1/fxATnpmp/09MxsaQqI4B4CJIbq1Q0oWS
sQ0GA3A5DtvHZQ1k6vHbmDeTIzYMjxulvXxDX8plmfMurh3/ufmePrYcIvBhUZLyeq+Ueu69RSh2
dIfZktjxwW9fBTzwhJvZ4JcD5WTybBKr8sx5DAvGeSQrfO54f8VczT55iKELNlmbmAo2KA8YCh4d
8ThijAGTk9dJfWc8UVXeMZqzgJRX9DK2/YJYGOWUITPDWvN19OK/cSGRH8BOxBhZeW8ike7KizgG
8lH+80ZWGpPJidGn3ZkC5Ek4m1ZR/GGLOWcB/yFaD+F+8ySEMKVVoRQ+ZyJUPdvZS6u7doTxOVYW
eMPSwKE3W/ia22LLUsJIlFvY9AdcEXbIcJv8QHONg25Y8c1TPE7kEifJrzU6M73jZYBS/3isSo7V
serlbRnzZNdHm8QN7U/VxKRmI88KZl72kK1ANKEqbprolrEd+o9dvN3PGTugscnobAYd2Cbnxmcy
a+lcYGk3Nhu5ob0ghoxaTccz8PGhvkAk5M9SxQKmJgNirFxfsqEZru6J2lht/J9+vMn+pMkKiDxa
5NjOW+ttIS/5GnFCjSiiW4hOm4DwZF5mBPXyXkdLphFzqdF+kuVbUlzGQmHlftjw/LtziQSCu2ti
oT167gPj66gJyhDW8ZuXLFsNrtbIvW0sYEelOLrK7/7NvbHCJgZTKuSeoWjuug+ySSO+U5ejxDGX
J3Y2kkiAD6ecohCxLoeb3opERLlTCwpTEf3ASgSELki6+Ya11X97xrsOLTzWyJfPV590wror3cPL
OwVI2gjE3+9085M156chJxeWc77lNqmypjzzmWK4w1U812JSqMT8JTRaJeQBVrB7ygeHudZ9CHFu
hjzGj2DufTQ0/iYLybtLxNCj5Qo09jWDba5xs2R8yrCTxdeiQ5jWCTpYPPpQJLjxsCkVWgX/JuKY
zXc8Enbr6saGF2tML45dZR5WS4xA1iPbMWneRaNk7I7yN2ivVCxCymLnOiJQ8h6yy9pq/c1UK+s+
DA8SmkVG8p5wamJEXirqaz5N/6WWcE9Jxhp8POLY6Mr5sO9tD1fj0DP+7UuIfb1CQpUDF0rMTncy
btCn5NmGicMLnMLUDdbdXOxjkBoQc8lCe2Cdu7BPBS4s2hZ3YhSc8OQyO+Ne8UYWuIHPbn3LJISi
isLZFzV+QeGkB3xwPPNIxr9oq35CJbNGRsLSLgJKaNNMHVBQI0n6v2z8PE6CTyQkjbyP/wAS19rZ
RzhNvrlKdOg4rzeIfitc4jFYYaW022XTb37QLSMK++vLCCIt3QB/25l5pZd65W1RyaQjWFiDgmIX
EssEr6pL9BA3qDGFJnHj/75kvLZkDFgIsKKa2oC0qx0zD75mOfgH9H/8vCexYSZPUgkEGxRcxBOc
rqzpNDfBDxxjkwaJN1po+sPn3nyzVAdSoOIRWzGV7/YsW3c2Lub82FLw8LW8dsQUbDlV6vW33MhB
tWRDyqYJ/g2sl/+aDGqTxrhRyw/wPl1BvA4o5TgU0z7dkn4FotekeDlhu2O53sZkP8YIl0eTlGEd
zMi0Sa5/LvUbm84UN2JqZ4Hwu2okXq85wk03Z6Qnjw1bcsm/q4sDE/BqkdLvll9BL8CBISjYjyUi
mMREXPQz3nDOgw792JA31kXmeX7jtRqK9PeVSmk5U7Mcgtn0QJvBKA78eJ36KFU908k4SKfg950t
L9hHjvACoENC2diSgUGz21X2XP9kx9RkqSmGYXFOstPk8w8v45sqGnkeeNh+LXibzJcFn8tBGxQz
JXIK2pcRDmlC5vJt/d1vLE2HFp57A3TOYyMvWREvSO3y/CN2IBhjHopxDUX0NgBZTUaECC98Nqd8
3EkjAlpa/QaaeCgRSgjszIAe2418ZSwT4vALqEDjGYoXqH8n1OWQpwFu0GcVb7wmd27V9JKQaWjE
V8UybY0vbdxeZfi4gnLvTCUxsTaf30HPnisA8YPXkiuv9r0iOGNSOVpn2+5Cx/mEDC84/sIFGaTs
aVm+QfA9fejTUPyCcJ0Dpd4J1nPQR5ErPNdNLpN7iKPua+O5+0JanXEJmKVb0H/4ZW8nv2bp17uA
kjZReFb3Uaoc/qlifyPvfDTTyNyE/lfNVCfTZw8kcd781Cr7lWurze2S2mnWcv0sBpE4YLwH1BYz
NAHehdgEcmezfzTOq8U80lh0nHoapeAUkUsvHOYExtKbRtOF0QLJk4EKaz7tUeVb+aTvYJJtuJ/k
97Ct9XmXZHvD5ueKsVuuLvR//PJz+6BAqSTsWpdmF7vz7ZEn3fI2XAcGkm36BVzHyCf8IR5Mlxmq
UvnUuayNQh8YDEFvgNpf7AWmMzHcdCVpH8LhZmDwXS5hQNZtQxHtBiLUvtuHI6DKY6y2uyhZABd2
x8QWTzbPk2BJtqNjn/ulwxy1CIXiGxkoyeFZXL8pJpGedA/TxCSvETkI9SXUMgEeOvrEeTAQWQN0
38qUJMpH9ADMo0f30yGeJRHhkql6c/crWVWR8MiY9cWgZAfs373ZJfabhaxSeVPSwFKHEpXSqJPb
rj+REA1IgwPDHSDCnGoTX8rb0cuw6bENEVhtjoeUP2JpbkxJp3veR6J3Sbx8ipiJzuxri0lD8WR8
7VKZnEUC3M7GaGu6G5TD6ck4fXlfFzhedP9Wp0GOZmERlx/Q53pMGOEhdbH27AS0mZ3EvIOFANW3
otx8hniF4ZM2rqVCpeThqqinKjhYBkXJj1j35dO0CN0EWWSQePtqYLzALjDmyjt/5tF2tHMb7q5q
7lAsqxkKzv/a2NWzixJm0e7VV4WTDRWrNZzOi78is8eAo47YDraFtJVq8HBtOl3EjYiztDkw4r/D
MjrZ/6DF3Llis4CrupY3PU+LRXay3Az2RR4bIsZOQmAvOZQSDraYK612BEdDqRtu0GTg5h6Y5cuA
Rn49lf9+ks/okthSs1VNrcoD/b5Vq6FHFVD4Di3kzCzx15fyi9gmu7ECxdL8DDWsCjm2u/LXchXv
sP7zjqR6Ws9bOqyqarb5R2lR74ibEB3jGNGWaq+eKGd7FHPphmkc/HYDHntdTQh5Z0k95UEvEaji
hwWlJQkxTNxxOtwDqGvBmh66nDshJr1wrMh8Hxf68JBifeYj68C684yF8hklckaMDz+nobeyE/Ki
4E1ZwxbOivcd+RdvlSK8ZiAgaH+q74NKu2DMUyOd+5r9ruAsC7i0uiHaYLOiUYRpR5ZOcj4d1+24
YueX+jUrqqaET2KPWUPXtRlgKP2i7Eh8t7zCcRiR148UfA84O5S0Gi1LMLevLzUA6CtTXCf8N0VF
t2l2D1YfiUK8oUfSnfpzxDgOl72kyh2+pKQh56xzOHVnhtvvlwlm8GjIOkXD54TYDL+4HIxxxTvw
NjQkzZVlrvk5YUVxiTU7gDbsQL1D5sSLLSTTn25sdsy0jJxrz6hFIPQAkhIjhSeHD+kAOaeiXisH
ASMTw5RsiI2S47gupgKSd5SWCFMEFvoKO3aePevw8pzD1kcA7MQAl4mKmVvcN42G8C3UdhYm241i
SMl6WGAUtUzeCeXEiCKsJJk1sxQFAPBscmRGG4v2MmVxreSlvC0gt2g7k1p24e7BhjRXKTkX1tmJ
Rbw6I2D32m2M+dbyYDeEE4ZOozrsSthDFSmm3Hy+FngU5b/5sGVozHRiovu4JBazYgiMxhk2ZgRY
+Dr0eT8XrRylLe0Lk2cbuV0xcNfMabeKzIKERBo9rLJVrv81+CVsbE+EgAHWqOhHkajnTmF9I7yF
KzOHhOaJF9YKoQCwUd3V675d5SiLINJQKLHzg3+MHmSkoYBZbAQis2lqmADNmItmTXixcxw9QwG0
OhQcKE+4smjH4HzFPDyrYsZiGnDFZqfZ1W7EypiY5iMm0OoeT49Y2I7RXiSL50KuUqaIxE/LEG/4
77aEMP/rf3Q7QD2ulTC5NbHqdkmtC1JTg7xnk2j7PBRmzXfmuE5CeO8agM9rdSDoa6O3oXVqZV39
tSAK+5rDisXDjewmOUlZpijjBAkLewA+l2Hk/Sn7REcbRG5+dpWBYXSkcu38C/+A9VU6tn1lre3h
mmYI7liYc18SoSM/geQpwdSxVeknH869m89Z9uXQ3igzXVOKvN3YSyzyD/XnWt6cTOjPO1p5jfgN
Krfni3rO8lj38ArTh+s3sI91K/0cngiD6GC+QOhnPL52CqoiLQPbCGpEdLPtJos0EHhSJ8DVZbCQ
ORy4oDGC6EAkqDBntdjbPoqSTIdXgjAhuMzQjAFKqiKBR+zHtdlFMzJqVuavetUXZ2yx0THOqqfT
esTiq2cWcZD5agG0nvTvUNGqvTfZj3H9I+yf+DrmFsj5XtZfw7hNP6Sm+JgNcrOzG/056XYLJbSa
x8NwRFoa2vnB7u2e+WnIqkgNnLZipwRqcqFuuTPWRbSqkB2DBSo9tgLNTWZ3inhlg6RcizOXrJAS
BPE4lJa52C5YU1cf8tV8Ma3gFuPJL+o58zjzEgE36pE/YpIwEepPy33vSzUh6qCbwYsevHURXs+0
1CI9ZyAqppwAcXzyjZ8sJiyxyd+Pj2Qn2mRxDJCvvM+/cMmOIqDbnausPlQd92c465CJlc3A52Ww
op6pv7qvmJdMseGhKjZZxc9Qzbo7RB8H2FbT+qCmmwFw/lIo+oihd8ds8clB2rRzC/wpCtF2/M+t
TWBQy0IdLQ11HJuwwvcKRWnVvnXz9CIjit19efh7q4DEmPSp6SyQ83u1Qyt56u1qUw0zgZzt/415
7zm26zIK/PNTY94LLDP6daIG3T11wCKgdZBvz1E/EeHDvUmXGHfh26YoVF/GbARj4DExG80Y0+s2
qxfBkonI9YxUJ/bHbSaP1iB1U6yJCy9+0LdgiZ4OWNU1my2CeSJkcFVMqiwEsSI7EMppvVaKAttA
fXQetq0SPI0RnniZF9BqnLevJ7+l8YZo5P9JI1PUR6p3R5rI0S4emf37KRmtf73O7wZv+w//vT7N
NAuHORwqi/BHFsc8k2nDfEoSH2I8uMUvoNd1KV6nHW8JdOPS5UxLxYy/+meTt0G60DAaeJY29pAF
mmRU9Ux32uhDKczD/iJa4UqP5NXV6NkLUfeDw1da+RS9OQn5Z3W8uYxL6aM78V9sjFdNT6dEpNY0
Gl1HFqYgkZ2n69bOYnYFMsT7gLUA6wCcuWV0ye4dqb0IYJ3AXgI0ModzodJjedMX3bRZosBAfjmZ
GkzQEBDkc5gA1WMIQIlOD5WzEN7phkXiuEXyD2w507rXDTjg2SwwNLWOY4pu2iF7vCiKZXYuDB9n
hzskKV0xFuUmNpw2EFNI2HF87v4Z7M0ZlRznqjRtssKn+ajVpYDaY98m75UIbuGETMiuCYN2l5OA
w8auqncXyAHqbv3gKHiXuX4K+7ZBo4Bgd7BqMZtOfPV4Q17r5IjRrfyps/GO907a6fNKPgQqVycn
WWbSfA4PmAaX8aXBC7BMrJWh1mlXxuJTUmrWxLD5+UYdkSXOLlZ0rHfC2iUZcF5ySu2PJN0l5Tzk
3p+Xr5jtth77kAclqf0QktAi5bAX94KkqYR05ZUWrWGgslXosHW5obSp6Z3UjKgVnZ1AfnCZHvQR
8HMoxYr+7Df/BaaYpF2qtGimhV8WlNjqP2rCY/jnYCoJjK2h7vHH988f3u0Anl/zTx2sZtAcY4cR
3uBjcMnxCGNyo2r4XeXB708uQx0mbzDYlKgZSa9d4TIPUo/8LZKPnSwUof03ouwRcfa9zbK6o5eJ
R8eL6iQ8WvsiQSCxsArOME3Pht+JnJi2yTr1xn/hCnME2NZ0MrKiHYB+DZJ15R/6FoJg8vG3Tph+
qVyM/FIHv/KC/CLbCZgtZ7Z1OL3zyMQqHue1NvkfMa8e/5I2BC3a+q7JkYQZ52WJ1/Sk741+A680
Z+gyI/Qblpo7EHJfRxjNMn+GTUtTX810mGADT85htUpCARbw6oM0fqUbHBdzDukvnT52BhM3SYfp
F9KuliziIc7FTnrffr4B8bap7Dt1mFf1dmeAx/+8DPtMgMOWkvVeqE12ymG3gt3jswks0OgoP61x
2sYzKZQsMGPuBmFTjNvjf30xgKYh/2tJYpc1l2gTfhxzRpQByDIX4RY56iuy6tViy9sj2fWcaFvp
7IcEMhA5VW+a59pMRO7HH+p21CUJDJW0Q7uOggTtxDTZqnI/+SnAAaBiSnXFkKWoiolM0skUqG3W
JAJ0MTc28KHH9ACH/Axz3u6pxr+UT32f0f+Y6uRSOSNDsQjVDSsjWCcezbgxvuEpA2tiMmwiD9aj
9K4JKKonqIrr70gvR57+Ps7f/vC6gsmH4xtd/X+9/xdfo0wlADIuezmBTyBxAJQbcxgJtW2xdrMt
F86wxj3xR4Z//kxDtTmHkdUOtdn6RFwG8FIqn992M1rTAeZvZByjG4flueVVtuktic6cQTAm18BZ
naQqchF1fHbMboIntiXgAIDrb2aGK174nCICHD5+3JQjVfCIgKRK6Cl8l715O5xauUkwINg6xGuB
0rqhFObP+Fva7FxeY7EvPbgBi+nkyYQjoAFJxAVl8AO85MzG/SA/WIXX1Dv8E5q0NfP5qO76zfDs
Op1MMv7nNqZs5pJMt894rpKV9xddPljjg03wTvb3tpD9jisN5SzBZcpsh2gqm67SbZSxgpCCiigK
dAypcZhPCZEtgd/Ri1iJJBvWTMTj3QKCrViFXY1hMn9kdmJpMs9F2XBSZ8yZUT4Km/JMi30mh/KB
eRBqrm+YmjLQN8r8DWVhgN5UPvprK5k1r2O/aK7SoEJeSvkBMkq7revtLKek7qz+njrmmjuRn9qD
S1o/EKeBPC5FXyNc3fmUbMZZlF6ej4srC3CRljSM664cAVL7lHfobzet+RXFPR93IKkUDvUwbRcX
0vTZfxMq2YdqAu6n1LqPAMKCbvsRGpxh9bujVtF1uFSMpf6i+XRQtQPG8yPhnlJ1Wckq1io0yXEP
Me23fiAUqo+2Xkirh+kQTB65MIzSdVhuc0jMhZMdtz7qp75VQg21ysVHZ/d+WbzYa4HeQQA3vGkw
06VN74eaeJx/LiPCklRIwCNVTeKe2PsE/Ma0D83sNcSToZ4DbBcCNAamuFg/ZBq3+qn9nGGiEmkY
a+AJDEAqlAonRrB4sjGfW7w2UHeAjNpjZ+3Q2yg96h02etWc1N9Kx5NZpJ4sgizkcezkSXtDeIPB
jOs9Mr3CGBNw1psONJ4rQTLlKFdGdXRZyjPfmPI5IZCKGZAwL2CraDp5/3AzfM/Hjyf/sdrPdgqE
ucQowZjqDsns9vEewrSAvHe6NpIOMB5pPJF9gv0+5DiG6Al31XAfj18ZbuEL7ugGRV7kyyJ5QIg4
16B6FfmOPixeQPUlz7Dk4jlSpKtWnPMLof20Opc7RDFWdM8urG1a+B6EP5q6XjO1nVCJBrBlviyf
KZl0xYpIRzWH0ho0TxQuLGD+PrzliHEYzcLcVI6rkJkbNVY9992y5RhJkOAKi2ytHpja9/xL0cJe
MYIL7Ki2CmMG13E3t4/BBb5cqD3sftzzLO6gQg6RGu/yVTNWrXMpWPWuJdX8vFJmnSk8xRxWuwl1
hTaYRpW33gWYXJICeqHfjzdfKxeojIn1p1HP7BqefuHkkQ6XFPijdL1wt4Z6Y4QOkT/KgZCXmS9P
C2hamWji961W7Hk+yt6iTAXnAksUvR+e5R4RwQNwfgxGx2ZWXu9PieuOyU7UDu0QAFEtyRm+ZMyz
ikkgxnUcmSJgc0MwzFy9eJZJESaSPU46bClsRtkJ9dpPR5oJltNJwcb3Q0PBAjZtjN4kSADkZXWa
JbHGHpgJ6BqDpwU22Ewp0C066A+WLaEHVZxB6m1mMDakWNG/DgONla0k8ako8aFZxfyRmggMxkoR
dzG6bqS1snrPpr7nLhp53URa4yR2UhqDWeC8AsRN/f3AzbZ6fDhntaAwpCAFFxd9I4fDdyTya53a
vh0fJbK+Auf63Lc1lsKDiCsNCvi+UENMgOGBLavW7qmbg8geIFxG1y+Tz7XQ5mnBpShWjf9NiKp5
5kVDkTAACdC3NS6yg+IbNTbe+KZ2ETvy4neW4QGZFDR/9UdEBGM4M4gWue5CZYVakdcshYbmixpH
886mALD3MEl13uJRAT9Q2tldvGWFd54A2G4hTttRKtSb34eGPqeNr3EdNjz91+Hw5A3C8D094aeB
PptwBcY8yE0KocxVeMI9LkM6S8CS2NtxY0B3ArejPCskIW8Gizvl0z6phaqLGtSjjHp0+ETEtfOh
sgkW/qgEphPt0UezEoaHDbWUZhjwBzh4k4k+3ibNEXxXNRS/Wselj3Pi/uvxZTcarCSqEWSS3BMU
9gI1dQ6L/88HBHFWQsY9b4YLWMzmptV9I6rmhenoEVmHcsczZPeTomiV3b/KGEdZOeYbwC3Gxibj
NW41lxETl6iLwKurYaSzqvuHKPEVaTVvPoxc/V9WHIcOFpC+/PG3a7IvTrcjExf/QDjJwUU09Qag
sld126VjlOh8jV9vQb//Oqm9oAMsThgEjaHEvBJdbM8w8+pces777IxhxNyeB/MxqNrnN+7iP8ve
9lF+mQNib7ZyTluBk8UdilEE18tehusPsCk0TznMo5+eAerbM3B0P6SI+E7jJzi81lZ0AAXriS1A
lLm+pZUZbkDd7Bu4I5os8l/G//BX2np7zkN8zfzIyhb2nuHhJriPtG/eS6MsnM5ZukLQx9Ixz/4C
CbCdxvUORoOzs72Ga3/p2aQqjX6B5haF1GezugqKWUxwiSg8qJC92pk77uJ72wtmaJh62u00hPDC
SSqPV/AsnFBUeQvBj7omO1zyxFK6OVhDqH+5ZoaPGfnNtHbeOaK9yeWbT8bbo9EO+BwkhqzG+r6d
62c4Jv40XNupbXi8mKFU9RtDn6slDAHZr3F0jjMUfVlqtHo1S2nrRVXQBmzdTbXMZheZ2bGdPSTo
8cjQGydNxNjR83HR7OcJc96a6f+4rSDw8SXnAqvVqkgC9IwZAdiRv141umQPrqLkdJKjIL526i0t
TY+y0ULUu7c0wYxMHR2UNZ/g7oDD2OPGp86lCdNw7y6DYNWgaGS3tHUPNTwQtGYa7xPGXtkFm7cB
QKNYoz57VrC6+22x9m40cTBii70UBVNI/YFCNzrrSKhUgArNwzb+ZdkDrES0n3WNMjJLblf3k1GH
xzGfVQ8yzqoOQfe88PcSK82OJUSo/zUOc2Sp26cMQ1B/qd7S1TpbFNA8QBIG3N/FilVieUgMX4Ye
bYCHLCFmBI5vtdy5L5v7rtLYm6Z88aeeszBBYOZlaaDHLOsqt4MTSKdPYFTs7li3bhELwYmBxJ1m
/htMTTQYIgM9LmhW5k6hY9SjJdyrYRXr0//kwPXFhc3YPjkzzRYBr/lPOf0Sis23AUP9Iu6ouqfS
w57vcsVlk4iCtsxE6+NP/TvUgHfEtvQrJNY3HDXf8mTldlVYZxfKx+zYEzVPrSR4JpyQVvZZF+LJ
eMyefzB7uccBzrGzX5XYmFfU8+azWx9bESmz/3e84XwklRlIxOEwg1Sw82roQMx0mfUY/1jeOmYM
PdCkeqPYQjSeLgZcvkByGE4N9HzRDDQmwxdufbUstNnPDyWxZ62JdpM+8AHMKaEOf/SRse49BEto
lHktgw2RzRBW+NG8EC12MLwK4fPuobQ9KArs0t3yfPn4kI9Q7S+PDBvgIWOGQL+IDYZ98o8WZQuy
egc8RtcZ4UnohzG+JB8tCFQ6dmaec9ZFHMFYnZllV60GmwNvXsGAkb/ZcqJGyZDjK1nDAnBuyUpf
yhuRJ0dHHws8i9gnV2jhdPdlwGkUHDKZ7c3w+MHnle806Iz+XKMwDbK24YumFu5o/5PaqyZ5Kx2Z
J0Dcw/BHPxDCZN1K3B0zjIng/tBupwMtww3I6hoH0VfPCpZJflGNmic/4VqAKqmB/IraYkfF6w00
fUbe4PpOdSDsElXsPxZEydFNdIVDwJsz65NWAAkRCWqciZMmx+Tc5lTBvEdh1z4SD5VhlJl7zO6i
CkjzD4LpxGgVlNvMagGNFdNJs2SQcw2wxdHTn5KrLTk23s+mC66KSW3aklG3sjUjLfxNdIC2AQfb
w7dADo0bcfzwkV+B6Ny/3h9Hu9Dm3sgRKfL0tKpSkhwBmBx8QyTxL5pTkuPjTv00NkFBrE1g8vK4
7FTZotf6g2SzxG+1wdra6QDJV6foNb3qiDOIwO28tNbLLPoOa4PPRiwZlY/SMVxny6ZxYYrWSN/n
BS1JBydJ2mbVo9xiLQICfu65RXTjso4XiBWvqFcJ8EHfno0310+DLe2RryOlCzd2533vY9kPGKfN
4m3hAFfDuXs2Gas13+C5MAwbM1PxbWrOFnw4ZNgJeSn/PF5pYZp5TB8djTfUwt/L7Ar9WO2JFpqt
vUQ6ku31aySWeTFxBBNG7mkfAJdjOFUJvQ+4oUXg8d4xbuLdIqJ2fa6RQWb9HR+TVa42oGUsF+LA
yhgLCVu39FdSB9RhC0gQsmDxLzoQdk9iJU5Vxzfy5cGISOlMd0hcdIpPHFHYGRGrTaRfZorYMEFk
Jsv+JGPSJLZBYaeJRTJMjCJg4G83Z5cvd9pr3dmxypa8vDsiIEWZhUDAXNSUEgdqJBsLkLd2SSr9
9JJrGpw8ieLsYJxUhjV+eyBZZqpnUuLbXTIg7F2MUq6m5aXgEPHhReFCb3byV4y0o+i9GQj1Iyyr
NOlMz5L6VcFqFZ6b+q9ZOQMfzm27+afWgAxYVJhguuyapcat7mVkQ2sU7RRFWUnLpR8zsc7Qod4e
/rV1LwXne4nHkoiiZojvyrA4lZfT1bIecpVpZothfBjI6aWP6tyxi3GUem9mnZUc6XwdqbN1GH1p
1xdyslvPfv7oy31TSi3qpjcUJ9wVA72gt8jQhO8lC66a2b0VwdEMwRzopXWH4FEwDex4tU0CXnhn
4p8jQxES9w4w82mhTDIk2VNyz0EEzhP19BA2CVfxZWD8KtKrVUJcHA80U2TraXUAt3Vns200UFNJ
sevSOCZGFFBLGYlLrKQsslzAAmFxqDe69yHc2d0NQEaJm2+flWkFU537pUsuKZHBRUFlCsSFvVby
TjmwKQwm9stRIK3c8bcyjriX2bKng4yUfhxr8fbgAezIyMd/Lw5bhm1lZW4D3c9HwgNQEgXG2HYl
hL66wSyUBmKbt4hR1iWQ3zZRUHxg6pCYjKRYu9Qz7+tqXlG1eAHoy7+WeL79WT59UlKYJ5ZGRDuZ
0ZNe/Mw5vWkl0YgDdBXcWGtQpjl/KICN7YPo1KygA/IZcn0quisCrtUcR4w0+MPRrAVBa6ajNYAR
e3MzaF+cso9b3fqysWDcz6Wef8Hhupj2hV9BrejPnPE0t9ZhnI72ZXsAHeMN7vOoT1HP416+6e8U
VFWGA9/02vCRwgCJiX/TCqqgqFkas9OpT6lL5ZxS4yd034oXSXMttwWfwUh09hewhe5PkXWvpyRJ
+PoFp1zkUGs8knvUBKw2fZt/UB8UKDXLhjsYhUXIJ+/cEKNip+rEfkWRsHGUVKgrD3g2sHyZFLb8
vpc8eXIyOuxS1nl4Cq77IP78PLUXLyhLEEpfN1ghJkmdT7St+mDwwLJwucNMHszEiUZm2Qo+BwjJ
30vERB9/OM9GlwwwbrK5kqNR1kewbdAAJf1Szj7wZVf5TLRieYABdLFEZFpTvd0FWLzb+zz4m/NU
uBag5aewV+X8I4cY5zTKdX9oPIVysooBU8zK3MBYBA3ArRSxndHCv08hxR8WkuF6sN8Jqx5VyQUF
m7YcJQljxOQ+/4ezoXqVuNLH4N3ZUGgOlW8a+basF77CHuza6Car49FUGx/3Nbf5rbgWI+25UrBr
AB9GVjLzjhKMHi0Fp0Gl6dtvBONpvh/yx+BmHO0Hj7pFHeM1lntaw0QSzoZmDUgOtakT2lmUbPaL
xb2lGGt4/45xuMHdW97x3ZVyjEh7tRyRz6c44ExDMLOfjC2cTV6qC0hDRF/D08pNER6HcC2aVJ9E
JYj+6jZdVRfjVL4L9hfqdjG1XDSxk6zHgWuQ3GM4Dt/DVO+bbn693wbUIMVpLQ5dL8kAjueD4S63
rupQksE7h3SfYkpTrU1TtKjkrz1olmkLcbVMC22HyS8wI5Wkeq1S6P6lyrDD1UNlcrGoX7NE57rP
uCdeVnYi7LO41roSood0RKldbU5YqCj+nXfLWI3f0oemhO3B1txvBt9e8sWdBQclaQm9DCRzXsY+
qRdRuGSckmT08TcUmxfTWvVC4OvYJONE7GJOPi81KKcDaF9UXzvMK9cPPP/W4mQ1CaSw5LZFpbYS
lWiPq5PdrHvpUqKBC/04i9rqAU3BPmDV6IJZSRxvn8ic5aeW5oupH5CU9xGpCrb7icJBf8bq3VOK
VZoA5HkmZY2EfPlymgv1pXIC65mKlSRe9VqbVZ3v2HEJoTiaP/GOq1S+IK3esafCcLa9W+DTJxaZ
Yki2rFSL/SvN4D7/dULCMLD5m9ZuInXwc/ir9zCUs7ww4XhWrzH94s7z+mMx3YUFvqRmWax64aWi
pK1bLKp5r1nUIjnsZfMX3nN0B26seDwcBzvNVZvZo3Mk7DfAX1FFM9bt3XBUnlW+bpthP/oYuyUy
dxaDt1JimwdMkZb6bIPjQQ1AUTLQJPAnrK40Dx7os2E4qR19NbZn4+JAC24cy9SFHe2NA8XdjdZb
Vtu6rZ82qyxr4YS7lZE6XyUAQ16tFJwssJgUmLMAHPNp1XOoa4DAyh3omajModu032cZl5naG+Mi
7MAZ8P9lHr0QvY05H6wxrs/GqgdXwm+a2ieiqO9CGTvwcsE/pDw1iiZXUYOyzADSW8sbHv7JrOZs
EOmDtP+f5ryu7AzdbAJXC7Z7W084eEfBHrz/k6tvexYizrDEej96gflxvGHrpn1/Ucq8iyVe3p4l
x3d8nLc0bZ0fVf9XCco94CFEGdLlrPOpZ2r+1bnqEMLqPh5KpYAO7uWEbN/ekC8EqXqMlwfXt4HQ
+nOvmVxtS/GflXMCxJN0Fq+vV/IgqMXt8Y2kQTRAIAkdRT0+LBrYbypjv8KC2FsNjS8kIn8Uiit9
7p3A6QBwytMSYFp9iDGzCSP4XAOH6PMmj2FCQwtTgBzrYqBc0dfXoBEFm1smfVtSX/pHZY8XCspr
bbbn5VOkBgUHWvkSZ9oQY8rQT3oHUMBQco0IfdZprA3fieyFlfOzbsfExWMveYHAif66pfDDUKUR
IqVIZqHNQmWlACQaj04qs3tG21O2Ddlbld7WlGvhsAF0zF/dGjmxAf7crrELNkGek9/YRJCSxqGS
BtoYKhPK2Mlg9b/V/MxQ/ek6rGOcHBrQ8Dx4D3R3jv/PwXr+cTVyKl0MeK5/im8K2GGvkI79yN4z
rvQg0Hb9yMUvI3NzZsubDa+Pv7l9a93Va1DQW7Wn8OsQe51FbhqccTds7qkHef2Ue1ntY2+1gGzL
W9L5LJSzzJ8yMUC4NxRPWBAwUxc+qiZZqJiSFyhJGpBQ8O0N5ilmp3wp+jSMers68udYexvxOa/4
8X65vV7ZvmogoxqNWFZJ16mq+9Waj6bbc05RE+ToOXfkLj61uQZmAkhsxavXYHTcRTRpYNpJCWa0
Z53Wj20wVMVtCRUS6F/Jl8zM1v7QApZEtbgQC1RnUuOnBd1h+HzS9WSv7bRXyo5JUlDloD+6GrM7
9zKrdZvtWrjrJZcCssgtQkK3fUpNPIzLk0besXlcmZgbxyb4vq/d0kHHbfa/ZUp+HvdneDK5/YQd
gqWYuHlp8fD5Wsdh+jTvJ4jCRf7o+l9sjO3WqVWeyJaVfaztIAmEMIkWTAWZdpn2XdGncUhvJwcv
UCC5vG1tWckeW9/4JLySd0e1Kmwn336zPXiiZZxdkIKvz8kSgkKXWo8ToO+17iOWvr1KqLvaAVHn
GiAZRk+WNu9GKD/txsJF2ngl7aCcx/VxSs2EjjkOKeRA0wZJag6yV/qQ75WpMMKe+HvgLoUz7UZD
YAF3mCowXBANPHJfJEcd1JyFk4dXMmTljDKKL1IMXmaWV4SD62XklHdI5AwB6eGqHzvy9WXckx73
wCz4+sqTNeHhCytr9KmsF3RGgoUnrdHJDIf5zNjk4Xwh/RQYVXsWzfEwjc8JF+ZGQCEGQ8rqeVn5
PLtsXD6DsUvAtM8QJrJBnvVBXRuijltob1UBDo0nbTi/XQfK9LtQmOXUrHQQ7fqBV+H2Gw/RMKMV
/TpiFg0K09rMMzo+aOJ2OhrPVfGwrIq9v2cR5dEtNMqm7lsDhZM/umcBbYIXQdne9ovT4GF3nyhn
3qqBuNmPKrnngxH+iK7duFClD2hX7fNuOVyH49heVzA1CroQGL4dhHvwp+Cas3e0F9OOR9tKimYu
f4b0UFRaY0z4Dvxlnj3GJUQSE6jo/2xPIAQ9sK04O5EzBUQc8q+n+GlR5UcJQCy5y3yCuZ95hC/R
N4FIT9vCq88LkTJ4ibx9/dzPDPlqRV62RG6nsEui6bgv0c8OT3S7hJKX7PvvHfzq4yfKKQdkmPPq
MxNU9+C2+pBU/r+3MBnfIsyCBmmreIameSDKeGgvpa7j/8W9D1pQgHx4iF3uoRf8WeVVTSECBGAC
cqZ5GJNI+L+a0Syz+AZtwMsb4+33P+vrQUkxNwxH/3RVd7HuKYskFGcOWwa+By1g47FIoIvOhrsC
3QtKDHYVu0Kp+a5uUaylZKtVCd5aGpQPxNilECp0yNK3I7pRLx9SBoZmEqnR9D1XbLmU+dkcm9DU
uCgm5jGj6DQ6YuZMKEEVZ5+Rg85NB+p05oMX1o4giN3u6XIZT1tKmARMAXTPla/Owho2IhqW0gS1
ObdH3RPKfMam6TWC30sw6MLwcrTnta3sucwzlx27K8Tl70BnKvpOt1rAqmxbTqGf1to8c7yVusmR
wgYTP8ta9i9HLP5ZGTHC6wkfnamQaRG3XafCb45VpqfY9EYeJyLySiTuw1E19CWEIwF0+kkgbeMn
hu3d90NFMeMs3U3VTuevjz/BNdm7BRa3rlAt4Tzu8sO/Ep8iJaO89dlejmBmE43ShVRYBpw9HTAj
menr5T44DZc0UfuLxirgnWArDt+/OUDz1m9yuBoAQLhn9xEhhHmZh4RbemuRU9X6AGzvCkoSWkOr
JqSJOjENn47aUeh879zAnME4eSQMNscUEh+T+fnhutRaZISCt00LH7XEgzjCgajYKW5yWuK+lv2I
tRm2jH7sp7IPj4TlWVec4XpqAamWOmuYP+WC+pDV+dDHDCdxMmIzAFfKMQApFwg5Ryq1jkMvovJU
IC/O8HT/97me8Lcf3WoTd3CEjUjkQ8G/Arcgg80XLa2lOxT8LafL5i79f8/XB7E1koTZi02XT79i
+sM65wLGGqnSY/URjhJZVjKF722zoz/EwABUySkk5TWq2IjVdBmM5GyFsl4bX/gg2866gVHPdUpC
oToveAZhHoUen7g57ZDzH5x5Ml3UHPUPRP5P+SGuseue9CsXUmrgLUBHbT2GfXyJjG+f+W0tDnbP
etjuBUBmul6SepCh0gYEj0plCfH8rWR00FIwad3INzQrMHxx72FBLeNRWwQ2jCJ73/CUnx97E99o
3Pu3fJYQPtH2m0ZBc8F7G3gq7iK3IPWLf/bH9GzvwwM3RXm7sJqBuyRWNz3CRrddJ9lPIsOkC13O
RAHx+gFG+1b9W+KEZUthkdzt9lJzRlauRbVwJrU6eaxcpvn6FgdLFU52kyVXfEchbxXnlo5Web7D
eUBNY1wd1zuMV4uHwnw133NHWfgPSn0UTV6kcUiB5D3bUlQ3ItlpsSmWWxDPl3VJc3SdQsB4TJza
ynF/4N6RJgO5XDvs4eJzLuwDegAZWtwOFlyIOqhnfmEJ5ipWvBIZnxCrATgjsGF8PAlxvS2x11r5
K2eoZ2NDlseiWsJcVdAHdbgvbNolh84fATlt4ZtWFjb1legfVo0+gY9EmiwAUfTuY5ryaG+IGufG
IMC5qfKLSIxNmirHB1HT/COt89coKryEBONUwx44r22N+WoDnCDHTFJkkd/fe9Qs6gcVeiD5Gjxi
7hyxTMxLNU5X2KzMMicNxQ2FhTvQeahZ2Ix+VEM6HXQpIFgjs6IKduYKjmU4NFrdUH1OimLe++ma
2DVnGEqpDqefvoDSRHE/BdGk2XBBy5vqW1hydr7Z5MkV72q/1FA+QmIZ6C9HXsq4SD0AdbAXLtLt
Pwy8zAbF/kQRGGCiKjr+hRCQAn22tQAztslbRZZFgsm64RZzAypj31KQrvFqj9yX3dvv9yQz/gsP
4ujlbGWK2nHgVOps9J2JLll8/u9uKYvRgUsv/YiG7izM/XACeWcL5WwAqF8Dt9TbitQZEu8XUrEE
Je94FUZVzYGBqnUDYnyNR67qwo99m/hGiXyfOtlOLlqduGv9H64Ly4sFMK9vk97IRvH/gTFk0GCn
2Hxj47oEiZ7+i6xw7EZbOy2T/di66Ef8JQV/FnJ8yzGwFXOY87GvrSW1r9lsHUa0E1TVbs9wGgQJ
okW3mBUolKQTJ1v005MS+P/zpqQVJzIDFZYHs79OD+JPQAhiDf56Jg532crnawNiN2Z9zdplGcP2
6VwzhRSARBq4GnHEQVE7I+z3iOQK9k0E5e8EGfxenIJ3BFNUVHbDVGEBiT0CTwHm+bND0nXvUVTY
qY7igZeABU371Jf2N6qGwLGdDLsXHhhjN1pCr7OKR5ikOATkHL7y/9oyak/dFrI9EdqBq5XqYLQC
ly9p8wFPlq9X8lpoX/0Xgl9NL9erY7gCg+GOULmyOxrfbxw8leHXKg89GOTfYaMdv8DJ+7Yy6iwH
qIceZ3zcKdRbgXhe4QwrTXlKNVQKGg8tOIQxBC6MpuYErKTKCxuC2y41Q3Q6CGyp4+5EGIT6oDyo
7JEgf9cIab0ouim7/yfuACJiYDZwiYhCqQYcEGl/l4enDZoe9eeD+q9znjK8rxkFnq3JNGvd58eM
Wk5KV9rn84VhwBOtMZfDam9A3hpt65/N495U1W97W3Yu4Sgd9oVH0a5M2CH8iHOh79+ruoPaKbfX
HUn2K7tfzwrpYNm0rJvS02EdheVQylfOkoyuuvbsSBaHqBcXLFN7+8wZ36WjdsRk70tAkIp7Ctgt
iowXWDQIO+s7/9kCuWCDTB9OO2Z6fQ3XBAvi6rtuAJEpVIam0ZPpglTNUrl7AxLO7CRalqtXrs2t
gVm7TYYhs7Clu6jiZ93RQoIZ60i9kuLyivi9kf3whqy0tD9jkVtTxBRFlBpXfIJXpsKolKN/LE/0
PheGi3+Z/ZE+IIB3JIv0SB72YJw2XXowA1hXWhSjSmmuu4nimPGD7rC4W7fKtFT6/pzrL4GQfSFd
04Nvf244Aniwhd0xLO9U+T3PErhzPdHRWvugu4Ou2FQ4ueqwOiez8kjQQMxy+cbyEitDddXGSj65
aHvg6XWfKMhyB/TaSdY9i6QH1bMjych7rPrTS1J7jEoGiPBkyBFW0XwpZNz3WAPN1K4GlNg9qYOQ
H2CJZYaTeLzDqzpzZdG5DVBu09S0cjVJD+p04UY30if91H8mJ9WqSWf7nnI8sAw1p0TdI+3GNofP
OVmSg2Agf4RS5u1E1rPujOdotaAflUpqAhsTmwZvW3lZKulQmyZ9N0HyQFNRETS/Sl7UPIX5C5fS
hkHVO4J2cl48n4wyRBNKf/KgXByXM4gENb39Q/wPa94PeyK2UDZF0zMRVAgvaGCfOvzog44f8GVJ
nLYZw4G5PXQZ4BYmS28p/xJB50FHlyaLNe0ug4mDfJjmsZnDztVD5iqv01jC19pPPBOsqas5ToQI
6Ic2uTNLvpnsKsESzPK46YZL9roB6rFhpeUcGuvHaMsoDqCEGH49ybbM0cEJdzdvyZ8XsPcuy8I6
eMFRo19SZKshBpPE2AEOjMuvzlFggtNt7YlE7PSz10RTGfW08rfgJQlbKfwAFf9GZjgJmrHtdles
vZ7n28qNmetkHIR4EBJ1jSZ022k8fg6JXn92IXM/nd8HEYMHh4AgRfcMMILUDm2bUuSgqyFVaHfL
naPr7hWFDmVFguNl2/jx8nH4l7wodR4ORjZP85RKWGhtPTZlERDwBtun0FCER9EQ5SVxEhVuzH5T
IyWlGx5z4Tlbhe9kyESWbKydhHz+tgtAgyB+hmQSLNk2rTV1FE7ZhXsW/2RQghUJsEYTSYJ1VcV6
3yu9ObzxMMB5thREuC4r2ozxH+qhLFviFyo8Hj/xwFp5l46lCCTBjrhtaAk5EO9cYrTuK2iNy+a5
wsbtEOhgVCnrH/LklKX/uhPEpzRs6qGwlwYtMabPt2ZaYLTCOhKtEuRarskVqmWcp+itq+IHGZ22
p8L+Nwv7B1r0t1A8zL3Xwbgn3hOggvccPb4oPJ+eNHmmDSLvJ9jZDZoPtl0xuMjOX7gBcghQUckW
Cj66v6tVTDpf/fLtKFjjtDb1Ttl5GQUXbI9kygEXZaUTs5N9O62VjCXGy5qoqbSPIeVqoxm4I2JB
JU1MNkrfKy/FuLwWLIP2Nx8hAWfA6W8lmJq0hu/TX6XJkGWXbdLzjENmJkNRQ5DXRgP+xLVP2ZJY
8gE+rL6QwwZVfxMT8bF5SbHsI/cuiDDVgeD65HOHo/LQ1sYe8WebybVpA8EDHEwO4re50bnBS/Ka
KQOuwWNz+LBUc0q252HAHucpoCYGbk8zFG5FtQegmzmAonEvsawS71aXz30Sp1F65lEsU/1JyHwJ
O+j4Mad7SdKCHm2VkTIZHtvuPq74de3bWdLlaXTrMBjPnUrs6TZuG+SnYTqzBy1ghjl0W9+CKk5B
E5IyUdoYqwKjKUNJh5nxwAzxgKgDKVanMaCZLdnp+2ouNGWxTc7udpk/TyVIFn5fY+OgrWmZoMHu
7xTCbDB/8wc0cXD31C5ylFcyyDB2lhRiWdMjxwHROzBvgrQSXHLMHURcFs4h/Hp290Dfdo7+vGRp
+Ftlj7wyTdWeTkBT2xiNQbuH6QwGzDba5GAjg6vtpOcTB/zB8WTNVZgdBG7Ofh1AB+e+fOW21l9P
AGyts+s9Xi2Ax3FztAd8yh1FsZZ4gcgbg3spr/DxPTD6D2oeeuALo9Fj8Kgvuz8oLZlaG4x/com+
3JnqybXG6dbPZw/JoLgez8POnOlUNZ9xNJ4XHQ1Qo2j2TwjUAR+KlpwHyfYDIJSoejUyWz4/AMY5
nIqL5qNF9HXLEpZKOlpo4uoMpC2YB7ek0WrSfM3YFiY09rflkWUNHOiAT1zfzWYNxyXV8GqgnNBh
NUWeUvepOzJOStof2CYattLgpIA2gg14xkGCFD2YbLa1iBB1/XnB0oBNyyTUVkdOQ6Wq8saPGoaX
gMKVd3UDRG4ZsTn276AC/Hnf/s0+9w1hifCE5yH36zaw4VLbrnxJWsXgqCzgg2FGJJBz9RT+SUU6
v4VZYx+Io69+2W1lHjb083Y3p2MsY6uP31d4v+RHaz2qZ4erjj7iOPpTD4xmN6NZL5yv4d/s6jTj
nqORVQ0SncHJX5FML3wn6A+hPRQKu4mKULC9gS4LuLlhGOJMaB+NdY/pl2wtt+m6taxuIHslMRqj
w+4x9F532pjPLwWpBO5QxGxvbeigMdwfBEnM+Z11umKlVUIWtwXDzsFSxeBNsQLd0/P0CKTnAmdJ
DR96O4MuldTwCDZaxlYa9nj5yOxBB6vqJCQN2J/6xOz4+qBFXePhB8xOFoGZ/fdOvU2JXX+YwYWr
QHuzJy88A7M7IU1ZIbZng7/slXHMBWvxV/VCvIPHsTYv4J5ci8lVMjIPocNcwUg+6N0VImjnugWV
gCNJHSYt5JtrAonlaNcNr0KbFT5dT6G6Jg/OEfZecj5dz9yASP98DIL1ir5zxisLsLeb/z3vXoJx
ksbmA95y/K5E1I8U/8kTQ8/8ukJ0xD7+ZPTqDuKXBEJN59nM25LyjAZbt0+FCZfBl7uj/zyRbxLX
seZIYFjy40sTodes6JcKLhz3Vv80ufrhLYU+SLTsi/4E0px1XL6GaVc8CQBkW2AnFQpRGbf7sYSV
NzNSZWhDIjXf1KUCLopjutoZzlmzC0QNlPwoCP8pRPh+vD7H6dt4xUg1LtaNSl/nsOcakHbi8bEl
vvnBFE4r9FzDqmh4KlUWStDVDj9/wBEn+SvuvHyOcqIaIvAZ8SkpHM7m5CNktGAAhr2mDgn7nGTb
NxXYxYfimNb2CxL89BpylpKsNCBgrRcHh/DWD6uok9AUBjfTbkcca7iU5mr7eoMe1iiSQJ7zekbf
t1ClKJ5I7MVsNK3u2r3kfJY54cIHjiUKxLrNFNBX5kcD78zF2hUyvdv4GrwKvjNrBJg5CjRqarpU
Eo2SQDVCFq784eItoccSfZTtmZiSCUgtjrebA/OaJfShUVTBqLFL6cB2M9umEaWypTtUDm00wdK1
Wp9tJ80cHAK7UAi7iFbMydYCw4PkzuUaN5YLSG2fLep+XdDAe5G1Bko+V3k62DPRgE4QLRekjmJr
b6QD4M+OLyslM4KxQlZlaAL8dkqnQ7Q/HB2R/BJaqPR+cnqSP3igl02W0qzAhWM38TSSPziG62b3
cOpCzwCTqAGaS0+AsRnbNRpy9OO073dCogQkA/JBJcAnwc3mJ/ZEnnd7poWbV4F0T7JX2HLvR6UQ
p8Ohrsr2+RTk1SzSBEd4W7O3NVi3b97JhCUydZlbPdxsBtzMk2He2ztWMeyBgS6hri4iILH7PUdK
AnwjHYjPQwHSTUDpAlx3P/6sM3Y0k0mgTfrbfX5TyZLN+PJIzVdc+Pd14DztFkZy9RWQxpx4QmgH
6dinSQWaoS0q/gS4nJ/K9ulIMJsO7ceMX2ske/zJuFSDhly709NyU3EeYnGejxd0h5CqFlpKyD56
S21PkgwtI7w4tfJbWh0zmsekMAV3VlbnVavFFpl3JzFsbyq63CIX4b4OiCk5Wf0NXpUyLgX5lcrb
rF4K+facwQMSHP6rJfgHQCFLkNvmRTsJIJXp2pJTMYT7Sb6uiRu3nFiPnufMx7jZL1OKzS9kbzNE
PJEfNMXVSI2QTH7q3fLj9MIWnyqlF8VCeCua/NjwMvH6jTWWoW0mf8ajLqkWcBAR8PaCKYtzge97
J964fxiTWFgx5gYTEkL5orBzLQXkoUfYeOjcvcwHryIdF9DhK7K2EW+8rnvJMUyi1slThcDrkn3x
2ldFLlVTHMc4FRot7WT3smu91iD+yTLVUediMhbgpCPFb0GVhV3B5v5bqJ8K2BDlyeRSHNMi3JBW
7uKhPLiFpD5GItgWMoOvsO4vtWEHtrQp88nXaxrflMV+QlgrqbML0e4koe5hrRppbeEq9DbjGrqh
Bdzk7UkdHnvokQ+hbJy+N7TuGZTEjlWlwNkyqfiKJRnIuvtGuUQ2xwC1Cb1vHdYFdB6prWVhxg86
zptVqE5XxlbcQ6+ptI7q7gJCZnJiuE0u1Y6Nc/oKBJR4xm5Vwej3mmWjltDUqXqCnZtTUUhAi+ZN
hoJ/RwF/wAaO3jfHRzTctMTj0CLzlNp9dq+TrOaCT8CPvxiy2XHWyGEtlkFx0/JjfCixhRS70E1z
u7AUvHRJfV21/8Ferpprn0DShKoBHTIT9JYMRSgGLHylacH2b+UCAf64k8e00YI+iRw3KAkpAFFI
vSDLFa0sLTi6lfEC2ttkelB6EP+xMN1SKcfG1mOGfOVloMRoNbOHzByS0nKesCfI+OQE82A5txEq
kU/tcViGTKYvHtw4hNMvq0iVLA/HXfXydxkbtA9hS3KcnZQudXOR+kjrBKCgoI/j9Xdgq/NdD6aY
/bue1ZzxXzjaR8YKOLrhycAc8jYjXjj1rPAt5wt7OhwbrxYw6yOzzthG485qjmyRWw58ztcbpvQO
d4LB5Owqr5zjJ9+Ar3ymdgGcxgu0xR9s8/CyIjdIwApvpTTkZ89a8nxadOanyvYMpqHixaGNAMWz
c+QrMzWkOL/8Q7ssZlQWoOXOLC/su590z9uTobVZQkmtjgFQUuH1o4aZKowiZfnxEAtLHd7vOCIO
l0al03DYzeFt2dtpLYCLpnfsA9U2MBovUJfE53fa0/1uGepHsili+Flus1cR/rhTy7v6P6yrolDm
wU3v7hXn4RXKyp6APkzv4ZS2yKmtCbvDOa2LQE5lqW9s86LySo2rLA68J++Mafcm99QBXShvqxwz
jPZTP12vtObj5U2fe/5wfM4fT+r18b/xqvmevbDH3QgIWkAheTQZry4MpWrXecWpvyrfVWGlUUb8
aPIWPcsiZLGiqRhKktwzQz7cZtqPd8hvZDbKjTACj3YmNsluDv0ujRZwS52jn1Keb74IuQu5I8Bl
XHYOAfz15Xxw+7RPys2Ud5bwECqE+SzParCjUF+zM3toKjIWtpQDof9DFhYynIZtBmB0nB9UaLT6
BwcrgqBgUIdFGJy7jE62I9pvPaueKzF7ioMLACivVuE5pCdyBwuRWPyUSLNUMRr/TwA8IGjT/MPM
dFCv0OGgdvkiWDyGbIla+UrUz4c9l2t7SdwBugL9oID85FCxRJMe9auWDBYwTkKvGH51ygn2Ze/u
yE/DC6bBMmgLhOf3TePfOBJ3/gRpYzAF8KiRH5H3XCdKqHDkAgdNAf5QMitaKv3ITGfU9FnuIyf2
aTCzuIPJk9X7cWBuuZxvWgd42kJ6xiyfT+/2MbZOJMQ2ElRg1GRvTdcI4yCI9QVocM0F4O/+MBHQ
pKx2ooIIEaxQ+TG9vJY+EP2msc7scz6gdgZzLO5zWts68hcraG53eIUilVDdTly/AjEZl1wcQurd
+HII7YUYZRTkSjZ+aNe9hKbpqAmxh2r49OhhKI4FKuVDSl4B3EYWrbdeV65V9YHAYDXbpHN7YHS7
OcmxLhM/tWKYex2ZjgufzdunpxIraVJQ00hpvHf0U83V866lrKbE81ooQ8W/oNEmhXBwp75q7oGd
IyJrFJuFcOW6SJ6xv66f1L4i47Q3gxKBiLZIuKGSMD0KYOhjydDBkNvoU9srZD/OwTSz81tGm4Yt
7HEcQfcIQInxVREQIuayh9ph1iauwE1qyvYZo8SSgW0VXuikKQxh6Q0cQ8ggCyCLy9fQo4KnZomu
u1xSDsOj5efbz82FxpCoQ78Bt1dLGJqStZxXmw5NZwK3mqee1XPMuqUF9sRMv8u7C7rtD/QUIwrn
MwqjpbGD3WWqPo0cbEz1lAsWK06cbn9wQbP4YrmV4OdXSnGE4VEo7u8tIPIltuAwyDp8atWQVDvr
RaDPId4AuDG5H8JYyy8DM+lvBzroYXZ+dbx9H1DogIlzE8gc1IcluoLkt5inCAly6cshm4KZk30D
sWBVhnyEzMvT4pSgIRvl44+YPwcKsmm3sLli91ZDsU0EbRd0F8qxwJP3rUNpLgG5+2JjiJwj6y+0
kjHDJgAWuMbm/l2+BQ9QhmiQmHseEGspj91kUtCRLG8M4hjURwTjEcU26SezvlSWzxs7hm0OIkyc
icGooLFL2rxAVBT/SHblUH7ywsZVNdqFlD+PGus2rc7/tuT8CXY8rFDe2SehVjNicDAPUsYRQf7V
4VqnAoiAiAhXbvSxYAHWDsbLb1W/izN0GzjEHmNOFEzS+y5S4fSJIt3D5HXVI0UHMWX1IVMw4zUV
V/QkHYbBZNp+rhXx9+JAh61HndqdX2oaNTETAmsb51/5qhcO5smqXmYuNE1755KlIpe2+RmFeALV
OpDTg0XWuWTaYgA46E38HJS8nQ0jL6aXkl5CP3bYTUkZai1uFWvzzcgm7tGlxdAqQTAOTKCKO3gm
qzWy65veLqd/hMjBF9Ln7hOzk/bP8YbKfszUGufV/Fx0qx9hJEqXuC26jvEOwNWPSW6R6hq1nUSB
rgQqQ7Z37Z+rgxStqLGnXmzQT4vjRXt8oebKW0juvv+o2l3f1N20KynSy1xX8OZTZ+oZWis2kfn7
Kz8YG1VDTSnAwactDZ3grd4EJSnmtXbPwsnaDfjgROhRhucnktpLQGVVsSzQZAqA1/bpW8qZ+KfD
U7nSR+My/GByasqXSrwD6mnAjoJ3hywfOhree3NyJgo6ZI/4Cpne0Z+R+1w3iXYKyMPU5F56nqtP
K/pqAdICD0tJ3XhpuVwk+0XXgtOKsdzyZgTJxZEIp/hqVUnQm8rMqNk/6I6nJ8CNlwYJUUOXQFTq
b+rAYeoeAbmHmZPiSpmiehYsfZRQV7MiD4m7xFmestSLGE6WR7u0pSJfAmcnSJxirvt4qxabc3ay
P3cGzXUlB7HeuBuhDBHVi2LuGDENiUcrMwBwX2yNjY+F2OdFhxmPBv4XTVTXDbrIf7f2jKi7NOkf
zIPzOb0RZwv4lrJNW2mzp+8AjXDRrgIkxz2ZmADAxfkBWPF4qsKofbQx0hzX1by7eRdEThoSKTvA
FPDErwfppzVPgMBhdploioNxmu/J+V4l2sEwoOPn+nfW7wrg0gqR5tvIJVw0J2YeFRzwdyO5g0G2
q5WKTfLUTU2DCX5GCrFpUsmgVNW+56pNRyz7lPCyI0obcCI80nC/MlZfuMYudVLe5FR+79AhCZsC
jutttX1eZzSb351Ho/V3bOtuxHiHXuedP4ntLyZFvqpmTeuuGVA0gg7oupKqYWS7hPE8MjRxJCvD
4YZo01ebtYJ4Gf4mTYwTlruyaMJcEysoxAwXSLo0gA1uBPQDtEkL3x9kq9duzbD0ybaSpU0VSoKn
S9LMaIoQSL1veHHaNxYOJeSA6hEIBGe925nq2r5UihvXQCi3QOGgbDzlpBG8yHGGlf3eHuRfvvE+
ffAsrt43HxxTDAmOKBMOI3k/WV38+LG2jq2GGTzHoTixFtVvCScX1Noer1I5TnSqgYmqz0WZPta6
qGXmb1J5Cvcf8oBFi4719uSDB+ulwvLqZ8eDY3zvh47Nv6qoQMScui00ek/+nxfz0zVU38oZj2A1
d0SrxdgyIHVhFtnkmwKGlshc8YT2Ja5l5vSdOvfzVEpEDAncHrbMRN/dmpsQEbS5g1gFR7wgEYVS
ss00St6+rpvbmd7AvsFwehc0+87pTDPPisCqc7dYyLT3TdCFPXoA4ViOexHjWYoxtfQzfSZiWKuh
4/7XgW9lbbLcYj59NwaoOB2mzdUPdii24Y6n9W+RrdW8L1lYqXISMxKvB7ogENqq2S1yxrQ2Cg4O
NJax6dhuoUmFaFZquR35REtomWGA/CkWZEYsRUAegJMLnf49wviQR+RX7vDYCTM3QCgm/2uZDBr2
tHwKXhEaEZ1KGN9HAINHwU8DR/XV6PiKj0Gzi4t+M7XNGUlPbcgbetxtpRQtwJ/X590a8GsvPjh1
esVQMDm6r9yWBTECH+h2+4LBhm46e+vYZEmxpi/79Slfg6lwOZUiabYXdThffZykixj/GCKYOoNu
wD/D0tItF1qoex8xDm8qS/+AoBOQ+1Nr4ULKrwOkt3V8yjgpMr5V/k+3udS8ON6i9omyQWtgiHIZ
SRmu5alDOiagXX26GYFp4Q1TJXtwUGLkUSv4hwXCmpaK+FJetsuJWXpUtWQoopHWp4O7z1MH/2Wr
nmVf29cvDF5NTCVJM3MLUPKislQ9w5MKwVOptT/rEy2+NCkdGLfKRriNJIbWRmLL53PJV1Cc65oY
oUFctdB+I8+z/TkEU7kRrBfpfo+cRlJV6rLKx3eE9J7xAIVq5SGc9gTUHrxUrhJrLidiEuYo8f44
GHKmrmhawCzaPe6z+zpKDnZ9sgBHwtNxHs3Bo+GvcKp/BcrPThrq/p4QEVO3P7bhJt/4m+U5nUip
BxARJon6ph8I5wKWs6q4qpHVVHRU6bSJTxpng0ZQapBoj2I5O1Hx6MiLtlgLwWtPE4wIlyaNQgWk
h8kxWDI5Wm7m33BFrgkilTKXGR0DAvOWFMfsF3Dv04SMK6dQsMDOcKp+nTE29Xz2byb795HfqkhE
Wi+wcM9nhZM3bml8VG6mJQTaSd5s+CmscL8Uah2GSSYSewW8a02OV0QwTM0lshJBW0RnICfXt0oY
d8Wx3QRycDuHVRBc2Tg1rvJoPO3tZUf3zrd71vvBZT0zoYHnReYdXNTLmQScigIDJsHCItZZvZs1
mbVydW6r8fYRgbw3pl0Jmj6o9DEHuDZ66fYOLXXgXKsuU3ufjdprwkYXOiaBgVYwFYVo9i3GYCVY
+j0Xs+CivpIpm3v7sPUrOmW5GR5cPwoy0xDs5WcaQXUZUseOGcftNcAzWNo9ZISZHtJKsR3qLO+Q
/aDWX4Q0eEfamY1KxOWFOj3toMVL/PLrdNCMq5fDeRD7Oe61yMfLQAAZx15eLLFvVR+fiXzsmBdA
y9wcq1o7b5FXtb7ByKdAycVYMmQAu/+wfExLAyvLzeH0CuFUdp7hN/nkRwkg+HWtZNqIbE2WnBZt
hnUgGyXyqogAORbmT8wY050v+gJE5WnbMIyO+D7NRQ5V+HsmNs8rMvON6bwnrSV66XinXj/TEfsJ
zfXRRWHlCPOE+cInwMAEvTx4CihPJMJvPT7yuOAoxM5XOQ1FjZqpbwlyxFLLSofM6L/OWnlmVrX3
ZFN4DXw4guYL7OH/RcrH/mGjEalkrVw140csfh0WcrNX1txz2Ubrqbbcrx4Rs75VuczfcqijaDiN
TmygEXZvNteeAfRasP0V55uBQVIOF1TPuI63IztvRin6SHiYjiPOhd0CUikftWCQAMsUGbR8m2T+
hwcWwidT6WhkvcbF5/94DJI3uOlvsGtIOR18gsnHxDg9rLEHbkum4FQVmcNUStBk4v6KCLzKkx7G
2gGsetTBpoNJh0BQeR8z3vlTnfi8lAZRGmrxk1VE0wy678Uhrgwjjfm0HxEZF1bWaGW0pxV6ezt4
QyMca+srReLpdrREiKP/Njpec5+rdkVwUM121aqIJzO9aFGFMA1Vn6QVmOqG9MoGPyQ4gw3cKH6r
ICyi8NXdjyjNXsPZ9nezloQnIIPdZIMxltV4H1UnA3Bpw6Z6ID0nzbjzo71R3i0pszpYRj1EF54E
EU5VJ574hQtb4LFTLOyfEcA6zMFqJoiF9gpOrj+qZDwg8eXtnNMRkP9NRDnZqZh5heQPUZXj6T6b
+lKCrMILq8I+fMIzGuOlOx1T3e0xzOfPYKdtnCNsm4FPIPhXzyrTjdLcKL/2lKaVZJyYKkpwE/tp
rq+lIWrw7jIdU3TH2Lom+Ed6zb50Aa90E+9jc0oEEXeXR98Wfn5T7pHn7JqnrQAcYTOBNIcL1CBl
NfOm/ap9Hh///gfEKXwb5ziVTaxMB2lyZ+xxjFnAd+hr7q7YWaukk4/5RtLxC4HsBokFTEvDhEcv
GVcylP/nJJbKkzCqJtE/l9XdRJ2t7B9aQ4n5SkbwDJCTtpK375DnO2pA+66DfyRLv+hFmswm1W0v
FKv9D2OYy4iVawNYJVBJpoYYQREtn0xkV0q7s7MDIxYdBKedpkYOUzn6TGGoX6K/cmeae+XkptJz
TKgeqMdGbDP3HusMYOxUrbTZo3iUfDqqraPfIkfTGwJ6slvU9VGQf5Ajyf+mw7ENp8cRESHUkNyT
Ju6NNMbazdIAsP093Mh6goqGKttbGKmrfo69enJEwBA1KHAdA228i4wZdJjaiM7tlzdDU4Fxul1+
V1yMjujbnHtI1XYZqYswiw9OahLlLMMT9cNK4S/VQQb1GXEgo2RRufHoXYs5UqncSS1qZ2HLy2Aa
GIQ9y/4EMUP3987YMlmDrzUlOUAE8LeF+ZUhYjjHl3CmFLRRPb3z09SX+JlXXU/vZBcmamMeX3D0
IBJuCkOBOFOBbTTvvcLzrmlPIPKsWoLGbo2N+tCsAdPfj2+P2rhzJXtLkHE1QLfjvdgEWyz7bsAR
zgOsjTwLqR7VPf9LPyaBUGQgEZbrVHDDAEYgyn2cV94/IyR+USu9MNr2O6Sr2muSZdHCBhcans6i
HhQCDf36/4QFOGsgpTat1lM6KfMyaCafAnjaf5DQzG/wB5aeOH1g8FKPqkJj3L/RuJTbeTQq8Wy5
f4+og9sQ4V9VHPB9NtH/7z4arWK8et1IUEkZY/RiA4FDBhAzx3Uulf5EGU++9l/lC8YUGpeXHgCk
NAmmrUe6ZpIJHiwi3onHHXE2v7LxdGiT0ke/W43quIn3KdOFKDGz6PsVwgQttsa91cSdD5hg3vGW
r0Hlf9OIYu0H+ejorx96nN1NUc8UYyEh2QSADctCAYf7ArKsiR3bS/kvKBs9puxXWzBTmLnGhqs6
GuFsWwdoUgj8f7TN/eEDkMcSYvE0zzHOoLufdD03cH43yQmJzahUn//HebVDcOmjutSIjbvhz9hI
Jf6PLIBYdVSia9LrijGVLnylBvv1YRBieDXDIYIyfGsZHe6JVSLGCY2bUl1Uqqtp7R1gMYo2AVhy
rPht9KG2n/mr4HYoNqoiuxue0KrmBf13djsLWAKUBF6yG6RXuZZre/loNij+0ITavCAuu4URAhjn
QxBDoj/pFLh+4sibutIyKRZT9UKSKsDRJxo9gJLHtOc1dm0ESmbwqVF2hzJ8VkwsysMdcIYNMahb
7xqv0u7I/1tkkF7vAoC//AtBDyS2MRonHGrx5Tbno4qeegMUW4Urg2AtDv2VmPYs8Z2arJhJapea
0CURD/FVU5URn2ay2AJJpqrA6WT09KjFguKi5eM1uuOF+hv+r7mzh9lIU/K/1aRszB+WOTkCT7dC
RSGPhm7Liu8Y7EB7chpN6JZSuegA+sLe20/S1okLuxrRylZuuX1dKmzfC6CjbVz62Lkc26xIcpu6
YwsS1PSEZplfhiIt5IC+sjVWQh6mnFYAd/Ujntw20UxfCMnOu1HNki+haPALB+Qd13WChiAGF4lD
le86M0uh62rXdCsGPs13mE+KW3mizTY2zlt1p5WYBHK4m5+ictILAw3Lf9OMpDT+TstlvmYbt5hw
4IsOy+KjLbC+qxlXjZfLGnxRx5iDMLyFdAg5+4f7hO9HjsS7XCngxo9jZHQMskKuhd3W7zLavAwH
6nEwVrShwuROExfhfr8nSSctqZY6UDIe0SqeshwLopJKckB9zOT/uW4sVBrl4xl4vmZGso4DKK4T
brah
`protect end_protected
