`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OH3qc9ByItKA4El3Ok9wxhDL99qXUCpp5V31QftcfYuT7dduDNvW1FLItAIbwrGc
QR09SiuSVNyEPmtxfUjICXwZgfua9pMGndnn/juN/M+LknW3r7z2qRXNPKOlhZma
HEkSDST0k+DphcBmdoYrIbIGZDCbZNmBbjJqTL1VU7g=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32384)
z+cQG8msDP0Z8nNJWMLoXtpO9yCwa3a266572n7FeDkDGEK32ZBvy69UgL0CTfyc
sjXUTYdMsmzMscq25joI01KWR5b0Nn8/yv1RoTlBwumu0fwcdHW09jPXA6bawPhv
PVvnEfBXPz48Em0kXl0vbPTsTXv5aQHKTe77lL6gf84itD0IGjnqneXC+P4fHtvO
H9jONNKaBAg7Ccy+2XUbi2KPpV5GrhnEj9136xeIbet2cG8Rywcd1UtsHHuv6NUa
Sx8RVq6lQ/2Px2Iopq4aIHr0fXn6OtII4EJ3/T6d3KuZemAXiln/6f1EDxaPzLjh
2K1IF/xDyQjpa4+lQy4WhFZiWONXdAKNGIaG3HfHPUSXOqubK9QBY/XS2ZdWc7xp
t5RwuqXmJkpDmzVZuIfR50uLvsd6BPtFsQJG7CRka070JEA8cAEBFRhzwN4c8x22
146YxDtzOxe099AGo/FA92NA9hM4zS84M70Z8GftiStEC98lF+DUjOd06Rnlse4G
MgPfzeWFKmbpGeYXf7VIKF5a1zaoOuX7AYyhxz2d0bypMfTrCYIBtVzXhhtpGDby
xKvV7VjXUCgKgZEzYSFsAz80/4Yew7ihMgZtFIdGxTuvVvCNcM5XWQKTE2ZxH2TD
3YCB4vWpQcplnV/b7Mmp7Hv5Js5+Mv5MTz4YjzvMqmTUIyTQcSRgR3nDICoBXojA
bEJEXHnNkKyJ/5J5yisp9JuT0Oihqqr4Z88XsJx1lcZ4BUKvM5IMNGNoHYSK7M9N
LWSJlpHu6dIGR+UajSuTUj1GKdFi2je5yTBH9KLhwdDUsXZtNGtZfUXHaDZ2aqvl
F/HNX2aa4dynS1iXNKT0/ZN7kIYpJv2zdkApV6CX/qYKVgBc8TWiViFtT7lSJZWi
0E+otKUSqVI17o62ihQHH0T+ooXaPPYaa0zW/di0tJQIprQtNyNRYiGA+13tjP7P
tOOoLV+6l1jxhAkm6AE5UxRn2P74twGJxU7N34NI7iFJrCEAb1hRYJpTH6eMuniv
q9j3hxeCVURXNpk6lXviyLYnVc+y0sjZeOCSK2UPVkITaNiowLGxANBjDe4mjsZF
aMZdky4bOUmLLQb/2HJGhjMI21gVuzS0e1iMIw8fN5XMDY63QdtnIyuL21VsBMtS
nwG37h3C6qRk+Y6iRe3sKtog7dbB2j3jdxHaop63xvu8zuRcNotnrdeCbzg1pb/U
Zj52FeDUacjTED+Rvwi3K5OekX/GfY9rRlQhZmX0FGl/kuP2Udcn9Tk+FNw/hfB0
TZNtBsSaulB1UZgLwUNXJDBav7zY3N7Qh7ePmYUQ8e+UpTV2/uqHrzcflAJIlJrh
NHZ2LSUUKoOCvfe54bSlHUN+7tl31oHn3bdUR6ZDJyFYFm9/kRu1VWrgAVakpECh
ZVedLeSgVVJen9zN/IYjgm7a8vxHVy5fmWfF5nq+srSyBRML5uoITPIA5muAG/9P
qtdjyrv7ZPPWtXPePwc/QKMLSllMhBf4zeA46rK58iSuD5LY7vNmaLNrTSU6IJ6F
yIdnxTfg3PFD12/E72fWVhYhsrkEuGgzQV5h8eiTjizXTySzH26Jx6W8LibOoAat
REknRgdRTHBS7Ah2UjvfRttmy+hsVMGlVjiR3gxrjtLMzkc1DUe6Ydm1OGCa/EWt
7v/46iG5Xd0guIGt2VUUQI0guWUIId2I9c47FsrTL4eXO4r6GsPyGvyFmISDINNn
+ceVYQhvzvejEKx2FI3Jubm7aJTVwYy+yluuPPhgHIQotc3uNHTTFEz1MIRCN0Gj
FnJGFAg5bTOQFZVe7X/Ltsk8G/Q9bZrslwvKFghx/Qvp4Q/GlFIoSCY617/PCLRT
fg4yd8NhVp6FNGFQ7Rx6yEpxKkd7y9m9/MHDsVr1LK4mn3GLcQAUbuJvo5GYlSap
R3bdVfCg2AwtclJ87sn+9JmeIfdvtYnx11XYgyfKR7Ciwis8Ud0FCR5LUdPbT295
0vkUmG/0Vw9zVhUyaMieaOCgsxTNjW2VG/a5muHwWH9NCcjfWJCJDQ3qXwTZ3vb0
Lv8jL/kYsc5KF0qFYXscybl7PceomWDqLz0mALIlDci0ntho/yzGxhCd5cuEc2Bs
k0Ks1PxkFSND39EMckwODlGOP0tuoB5qG/NH8Ur9f7cyWm7e4P+77+dFjN1+RWR0
V83iDOx4kr4hsMUbgMNQlR+co02lK0vi/JfNYCp9K7XR6w04/ytdAhquu2Nea9bx
DJ8sxxzZvjyRQ8T8emf1q8gpJ4IG8tTFiG6axqsbJ9y0+8x5C2tlxPOfzX/gS78z
TXzVafDWKtTltcVizT+kJ9a2SJzW2HmZuksuyj4PM90jLRTGdJBCgLYHaLBqDiYV
rIHPcbPKfb38KNFXgJ84Jwzjgt3ykUptwJakXPEtPo68SMoH/mNkvWQjYSCOLQ+k
sL8LDb66ICL2s+cS3jNjtUROWzbCgLT8QUFZJSIFug/EG1NpaJSiBTE4KYxpWuIH
0DwIPjpnZFCleOwnMv6jwi9s0bVp8gVtlQrDkeUCPBZGZn0Kuxj+PUF/cBt9bC0y
s+NY+6aAg7sWFkaV79gQdI02V0Fh/xRgsoOgumhZ19ZMc2uomn+H9zE9J3x+qY6Q
fAH3N49lu/ttsDxd0iWhGyjp68qCFVtB+jBJbSF5lCIkoA2a31JpKjNUoVdvyeMu
R8QzFjecS+tjJy9QBGNcPWTrp/uRr0XIczgYzN4PF6eOFPY8lSxPMnpcLXf6oVyV
O0qIgi2MUXsdrnGnXnBgPl8iXdO7rEVYLZTNp4WMMdW1x7gLS5WHnatV2wn1ZWPT
0wk2YYMeNQCvoPzTIZoIUDN1MTdq0Ox6cf0+OYXhUTEKemnt5PIDAroSPPeWB4Cc
Z5AjgBUGMjgC0az0gwa/dmHFzpjcRvdOLude5CG0E7qbGa10LqUntlv+hGLOqcaP
SUyNcmYYGGCRGHCv1stYrq5scTv+rgXFxifUVMhcC3HvErpYHJXjUVkO1c9N4FDO
rD2S+AQ4L4VZr7G9SMVmckFN/5q/F63YXxByFaosxDWpA6S44/QdJapqqcQa6Z3N
5OYWwQpjrz4hUtdCP5od8to8i/LhiadifEbx7lbABOdg11w4VYyvHXSJu8qNDPlu
ZnNleKrADwqaNLxc77TwbcLNx/aWo/wvn0VXQb5lT9CTmpaigt+59IsFZVH4uJ1I
BRdpCOn75+F2WyPL5qcfUeTaDOpkL4B/xmM5xViDWqjCOe2OSsVz9yyd4J/syBNu
I2xWZmoAXIJRphEyTAIYP2XEu8mdYmoi6jpSP+W8IwEiL701Z6BVMclkQ6yXeQLJ
S+kmkOj3gmgm3tJ4Z4Yaorp9p+Lzw1rCZF0LQhFmULFUbxGLy7C/44ZSA2RwCqdQ
BIsGOH0eoETfSkfUqPWDYqwrXvOqmkxWA+nt+OrqAvcaxVYiKoeFos+vLXDe7TlH
RfG/vLvPgCpAMCioN/9np9j9L8EWEuHiSObyIP0eHGA2oDlBzPuHCUJC2NG15vA/
NqK77pqpbNPOftvdr+aQauNnod4yNNnc1aSM/SCJczhXgXeWQMa17ISu452EWmLi
EIfm5W5C3LeFJEnTPwDAB/WQKw6rOWgK3tdYMv8bEBXfrIU5m7y6yRunryj4wfaL
Wa5c9I67IQl+sW7Q/tzNOm/28GIpPoREPmSj4pUZSBFwWIP3toJd9MbR3Hrmeg+O
3nLzf3q/38wMKxPnI37gAPILkBatMqthTfDE2wX3807lo/PU3YUzWSkYhQuJTihd
rP42KefBuCkwPIvDgAY007leiEED7i0qIyAHeqzjyAM66xej63maL4yR4ymrPl1g
2kv3vChBUlygRDqdtEWKA6NO0CoErnHHAgSIi8XgaCFhIQTtUGYsHmLe+ugZpMWm
exKbxb/hCaQG7f7M7DNnLfMqnhYnCmHeysPAkD+Lmh6td8groVyPdrL5iHUQ0WIy
vnHnIHvLH+1GxI3sXaXufzN4Tyeo5BuJpOXeQJk0OcUSisIs7OeVEfawMX7fP8yK
hLmRd/swgZCSz7oNrEd4TMeFGUqNgwZxkMCeYiCFdSWrvIq2JFOYsnGyEGlVonyK
//S2sYHM6+WhEgGbbek4wKHfHRynlcVi6+Kk2SL0pZ+EFr2G2wZ/feazZZzAun0X
8OvRhd3A74kfILD01tsIUGrZvZJSH7jUfrhK8QeuBnd4YjtzcjEOgHbSMD8YO5EN
EtxrcF8ZqXn8ColTgoC4velFSVxcn61cyMAIL3N6Ihm+jS5WjZuIcTnrnIKtPQBh
VbSdCO6U2L3+Z7NoKpZeyk1vFa5wnjRbDYApbVpLK1gtbe6y4TVBTACsKIbhmj0W
U9XNuw7vRNgZp4X2HAV5t8BzAJz2/zi06xnj2R5DujkwVem4S73H75rAs2eojZUR
1QQ3RvrVfAKVQg4nd3PVg+oFoei31daP48ZesOGdXU+RPV1XRSYa3v065Tywk8AW
ipVraWFgQJapTV6gwJac0aZF6qvp3bFeapAUrTrM1V3fD5FW+2KrudCzdr24JA7B
QjlGLdhomg7sHlWzJ536ehfFgirA4KZhix/nj5q/gN0s+1kLDnHPBLQiW+Keq0i2
aa9ML6NkxrPX1GQU5ro5dfEodvAJZtrgs/8efFrhCNcXM5y2TplVt2TpC3cgXtEk
VBKbIIkLwDyHl8Bt9q9bmZXWxNxMEG2Rs4POdJ0bZDJvNIB7FN5x5AXLlxf9EGM0
wSKCIjePZaEwaRqh5oWGTapYeAkGcjsmDIhvav/Qk65hwdGXWsyWwyIM6lzKjmnY
M+kDGe77jnVshUfDkfss4eJn+2uffYZZ7pbe6Ll69u0f+hUNFIhwOH35N7RybJIt
wQNnPtdOnukt1Z3IugNov19U42MpcBNNiUQQrFXX4Gih+lFKPb2c0hZz58TiJ6uf
qTaf8SYht5BJGLNs0+ij3wTIx/rUMdf7t9mAVXYIULj2bxifaOO587X5Q5ufCD6a
P20XihjLj6rFKXCIgzjvT37hhqM/0FvZ/dnSmwhDRKEFAla/aqGSGEj9LLj0/GM9
xLaNUgL8uKpACL6uMiKYHPKIrJTOW25FOIXIKoFp5fEFHXebGDP+lNqjsiCboKOv
iXaZbCtVQrSdtxq7uKm/QQfP6fdevZt9j5Leo3gT6SUtGrGhlXQcnDRNuFnQ+WSp
Aa+4sggVtyYzdJqZrrDu6TgfMmuaES9YO0OAzcZgsozdxsEoJ0z9yBnopBw08wIW
hGC22LmYmxUHlsw/2eRNfeMsbDuD43H12Q7AmskDUL9oSKHlzGsBvAbEKV5eAA0N
QSWDUHakd5PBZ3hk0n3dJy90UWtplYx+m+rKNfP29tE8O2SBSg/0bqM/Xzeid+zF
R9D+4fvmlLr3EmJAJYuN9wbNqJkeuhz/SizqLFRCjwahDAld3V+YPfRy2zsPD5e9
bwun/bA7WkTkttJjnVAt40Y9qr0iJkP1rC1ywL3ITZsk9coZfrwmgdB9dIXHTPtQ
txpOcmcXHAvLlujhi5cLHwlyDcpheZzScRlo4YyBSYNEyEBL12Yf+hAExm3zzKqn
dmgZCqeETpCkOI0tAFvShrq/Sk9R9Uf1eOLQGVicFch/Dn8mZzDix6KCMaIvfU3A
PpbXK9z9iFyyYJF25rFqgQl9z3ZHPRWw+6YlqoJVEcJQzpTQPvTSL4saYx2TGfLT
IlGzDFNo18AXqjNyEZhNL/hlSB4+DNuPeXkXcO0N00wTWF/9Gag4o2lB7aJaAcAt
do/z+bkHfdCPi74tMAAheusXYN0MXcrZ4Ho3OFTmYn0WbXldmCPM2PEaVNRHtADe
uVD5IWFAwtb4MBSPbIDu+2l22zxmoLK6VG0MVMzpQz+pj+w8+VLtU3EtMMB8Ddm6
dLWFwh5k9jTupb+5MGkoZ+BDOAM2nPwh1Tj8ZuO50W+6fuNEsekDokKco9X6W83a
tauD21AObCF1wiBAd/dIV+J1rhrSYzpKy3dGzUjrB5kcYVmo/YzaoCz30egR+CrV
iRg5jngABUtuhbZseQmdTtzTsZ5aZ7hnf7AgggOkI1S0Cawrqdi5bCf0miVTS77L
7W/fAtOJmZ4JijHMNtYtK/AXR08yFOWCqSRQFT15eaDkXHVAnkq7HMzOs0VKRXUO
rryX0oEQ4V9Bm4IC1oR/lYkZmWerOe9m32A0BOA1yC6FPYP8uR5+hw6YHDEIniZc
DY6FDbkTVs5Suv9qFRakfg0Q1s3rPASPEUvO0QQDlvteu09+qjhMD40S8rCS/bC/
Z2GE/nfB9z9IaNO0AZ6bTUB2qNNNQHNf+odt1WqUy3ItSF4qZzvjKteonJqIYnVA
lP9Ta8eRb3/6AdQhksO+gCQDxbfudTeeciYd1BIJVvbMseGip2whK+O8IZQa/XPf
n0ajDbxubxtHCDz8G4cOByIQYTvhf72/CtuSRt8ca6IpwkmOrNaxdVpNSj+A+4UW
9YPUdaho+TPS1FtRHq9qqp67912ICep+QVEeEUrpwdF89oTJ2YeoiowQAm7A0pqb
Keoey7jpk3bD/0yIK1lLtmAkyMe1yAtSdwB0g1QNTI6wrNwehDWPXxOV/TUc/2E2
mSHFplqFM6lB5lFkIwJps4faZpyw7zF3/zIAxlS2RaMY653O97dlIBND1g4U0lEo
DGkzM6y8w/WXdhDp54haP22i8faYibRSLehv0BcnznrRvGohbVO5YOahEr2P2VIX
Hd9K6lFiYnViXp+6YKNNZKJVFv/QTP18Bi7UiGjTyPUs3lh/aIkzOJXxWtfZL7Nt
qPD6V2DMZ+JUWdBW770jjE1PswawU+S8yfYO5eZ2f3GsOvqLWucyk87wsUJcY5qL
O7JBvCm9Ex9mgN6u+kRD6K9fu7on39UnA27ZF3ibD6W/xanlYKMt98GdkTMwJsS3
ePWBOnqfOGeE1XBkoKlTR3gV4tZtln3p5K1H6afh08K8D10oFENCBniGZESTiEyr
QjAurqd0v7rdCP7jwUASSKNsPn46BI5rGoW9eG2WB8a8HeB4VAWL2PlYWoj3SXdN
KnqpeJZKjjdvB05Tp5eSZGBTV9KTqZrhvfOsANLXqhe8XgG3+Wq1WWb3Dv9QnEij
FH4bgBls+6IBsjkL9rFYmh0AHq+YJGrlhFCCg+G8Rt1pXuhhFYUwTg6dESAUV1DL
F5fcrKtd+q86BjYAb/B5bjIWy2xCNFGNTaUi0yLkUO9Lno0ZyvhTc2ffYDd0yMBU
wvzi6bGjdyKD3xKrmNQDQSO3PS2Bopsi8043/aLEGcwAKK0GBdwZLiSNClqz+DlB
2giDRrbG4WgSR2ATxv5KxctQ6LaIwex68BhOdEUMEMg6RrsfndvHPH4iQsj62TgI
6wGmT41BAGRGRa6D4Om7Em8JJoAyNQErVT9B0a7bj60iEn/KjTa9OX7YPe8rsWD5
ozaftNQNxYwtQPllb+AAtJL8Y5lbDEffuXXtgw4FYWCNpGWVFdYAzVGh4OyzMFef
eGLNMl74+L+ewYm2q5iIMv/dnVYXfL3gGvAi0WHj5Md6bq8MeTyrxh3gU+rSaIkZ
p4DdYfJCv+cGwtGUv6c096lBaIXQip+LpW/RYVFgfsOCxm9i+nRueWPgHDY3YSAz
1iF7McPJzy2bopzoc7d9HX4DUm3L5fSkfdH7qgZnQlgO4oJoVgNboWsd6K7+wmKW
SlsgEXlODduR1Fjb472va0x0BJUUI58d/9xUOCs63sddcG7IFGuzTH7JgYOREqqR
X2XBrgoyRMjh3OQTKKGxpT5U9feSYgyE7qmMa+lBP9ojY9p7CIn9LJno5rOhVWUK
zTFFD8qQzKlkxnEvkLlYtkkN65Zv7TbxRwuogB95Erv5/35EvmQmjNRI/cEhCytL
sOSODAAFkoUY89DkDCSxaf7P9Ls5cq3gxKsNQtY+IHuxCiqOD9N7mtosFoy4U9Oy
ssJjkjNutpf+5Rdun8e5c6j/Gb6jhHPmWY5gQDGNO1iqyNGJy5o1JadwLNvqIAmX
29vvac1hf3g3ThhT+8dhHkxNcim5g16lRFaY9Hzarn9cga4NikoW0fL0KLDnfi5K
4cMC21ldlfs4/AeSBABQIWZrmU7qMdgNHQr0zXNHmKfwcJpC/1/opbmB/nmRYFVT
LMrNpzC41Eo1NNSvUQrhL2kSqzg4wM5fMIkJ7GAoa2ovJ4S6w/g0BFqESqxwVybM
sa4RkSAC1y5sviVwQCzsGoCqGLRHH5k5APjLjiwhoSykiduSh/5/yseUKzIz0w79
Ly3zzyYiedGCfij3OCubGfpsaYkdF8DOEsh7c7rpJffghdrOogiLtcwngo2Thsc6
1p+A0vSy3Lk67hIOnwyz8PgMN3k9G0q2F2bPJz2W+mwMfmb7mIEQG2VvdtRp4u39
G5QbzlxNHcL6/zL1VNUX5+pTGIosHYIvreFRdBvelBRFbQOb2bZ7kJl1fEh9mSJE
e5TYHnc/BA+KvNbX+g16lkQc390Zts1sSmA86OrtMmzB/gXX8P/PvFV6imlznG+L
4YBt2QyCUFHFQ2N5bctq2sYvmg0qBPdXZd8bWGV2C7mqYtoJEE1n2BK7dsPsYi9D
3P/Zjgm3a2DdmxEQl1Os+A2vibn5N3cdGOi02C6XCjG4mnDxLhhtR+GD18/ZVfp/
+LCOYRG4NIJMUCOeZZJO79V3X2c9y3K1qDANVqTq7e5gglEf5rDl3nG5rgiKeRW9
e0cQh78UAmm43nTPYbXsJvV9zy3MBxcRu4y8NEcN5BBwEauhffzVH7cOMycv0w45
8Zl4hd45XGox+OmWhM2pCCy+fuhdkItWrgPM/iacSq7WyHgbCzYLMPOfLAmX14Sm
9oAF+xhv95H/EuPmVRX845SMmd8lbMFUxRmAIgXeq0WxYeonPslMuBDCIyuE4ZcI
CDaGAxGlRJRc9D1z70JqWtHvl6iNmVMiyojjbqssFdool0u9UQ3QLHkKefCi/cYB
sPlJGyQpN7DZc87COzuGiu+eWCx0+tGeHxg8/XzJdRuS+peHJc7dcTyHrd3nJOx8
8iLcsx3Xzb4FXb2JL3RI27FR6z/arLBvKAtNv+pQB4tEgtUHAv43JsFHqJmIkEaY
8/08lNCR+37IC+SZo4JQWtFbZAUFEocZPsXsEgV5+anSUZXDrJRBfDJkH0Me6NNK
mMJxuyRnZz0o0FlNBtiziWi6lDcc+qwd+TKrag+XC1dgHfs9Y/PrGULUX1oeupHb
FRkMh+Th0eekHJk80AoVdcFUs9kZwGzT1iWrVXhawfR/ANapgeRXeoKQWZQlG6Tp
pL2rsMZM+K4D4dy4RgxPOGk9scWLjN3lct5+2w+XkqOdIkH/J6dnjUxfc5YW4Y3f
KpAQrUSQDWv0V97rh4LpOsnoYq2ukFQnlzcMMaJKqx5Cxp4uBradk+LwQg3MGvL8
YGtqXkNLSInxmdqJ2D8FYkByODFlcBGlEb0jSLGcmomIjxuVbHHONU9LDDjGp+vA
6sQ/LwZVgYYxJY6o64rOmWSeJ50G9dUyCElVulmTllpoNn/r1kwO4Zjwvx/Pxs5C
AHtQmt+AZAMOMzphZK3nmqzoJTu0BFzMRuGst07hR1IusfW4ohTI9MkQHX1m3aZz
DBVG9FNcedQhuinkfy6TLkp3Im46fBDNd0knwg19mvOtU6NV7BlGUSqiN5Kwc51I
NYcO/XBiawK6Fes1J6O781mxGnDqVKqn3OlQK8NSEO39H/ld8dRvFF0WVRCgZulY
nKdr8+1M7VR8+P73vyPap3C4YGMBAWUfcL91zSo/dB6LE3W7PHMt4uZmPgMjVsJH
B25lnhstTdpK7Gedf3ycSvS37LMsm9xkun6BiB/4MZTFfYG/61yoz6D0C9guhMdx
kof+LFqhmxhy955jj0OF3Y61UTPFMvd5ycsHCm+fe42kE/rJvUKm9cvu6hWW7pEU
HNd61E6rWY9UD4UIROeaaPpLsdswO/YS6svp/C9xXcLPqm514oQQbqaHzOnCCAUc
JZPPyBo3JE4FZ7V3kizkYcAq2HhdKkgc/JtH/pbRld1Uet3yrohbwkzk2qB4Ov7e
ch3Spha+9Mk/GbwKvCXDqDWDbwG1JOhU/a1Eepg9S3+V1YddDJaulf8lzBThiRY/
FDLI3fjFKKKkBN0sSMC0/IZXJW1eEs/ubGmiEZXnR3qA0xuJGWopYmLS0jqKMnEJ
c/bH6pbOMeyAgbEBXm0k7dvrdT3XmKefTNBEF0HEujJ91Ghs+ApDpdRjSXc8EUsL
+avFpYiO0DmNUHxa7Lp+as6TnlH0ZDYV38qHB6VAIUVRa+AsCNuIjMMP9Vkv6gqY
adN9fNBsIRnqpqP4VwpfHzfF9TEPVd9kPzK6CBm3sI+Un7gWBhDCTUey81vQcEp4
D5/1ilHMadqt8b4+/r9H9gVeBGrRr8ZEBiGSiK/PGv5FapANbKyoA1pMRB7iKYzx
VM3URbqHVJ8PPdBpR6EAc5I+jnjD8S9YrsCnS+ej6IeKuSZGWKXPx6B8AVfSvncT
BsdzCwpYnOARxE6lXKB/c0bZ+HN3MCBfbgJ6fCR7/SNSZh8cShiZFUzHJaNHouPY
K1+HVzmm3Ev+LVrYRiJhj4d5qr7jShtH1hpbFP5SLjqRmalR7OPQD7omGgn9FLfZ
/meR6H9v48Gdg0UkWBWelFRUMxjatTP/ovg4Nz1Xhniss3vC2yAzF45EyuZaIMBl
WmTVfF9C5JI18JiqUeaYRwwf8tUY04RLCS7Si8ZCMHJriwRTWH1souygc3sIEGPw
zk26LBsXjK/Wn4Q9qFpgcOuOSSBztbdKFrrHTovtxnlPrGrRyXI492aQNbn9CEGv
sf7kLCna65ANXtsJsFcIsREIBpIx5tXNZIqS01wxZWDVkY3fcyhyo8Q+6aUV3qZt
19ywBnpVG2umokwPgHGPJz2j8QD/Hs6y3qfEuaroAu7azJoTTHMA3O5Sh7lJ2Pso
5WtTloI0aQUcqwuC6hbRme/8TukGg+LzC01QKNd0oPGKm/PYLfATtSwoggO1MPSb
6r6D9usJZdaT5+rl1VQ+Y/9kMZkX4Rl1lOH6fac/1nnLheGd5wYTsoI6t6JZWqeF
ZxrcKuToHmT/VWCsWKQP6/tBvIY5rJgfyyPIF3cGOJwOyr4RRchnOPnQ4Xo+9HTP
4X0yAee3HSrGoeNNL0HgOZ+NnyTjKw4gd3wWB3zcuwqZHDw2oDh5wj26mAz/Dncp
crzPu7dasOfcwooQ/AQKuRmkRWM/0cedHMkW/Tv4o58JCETf6NkOgY2s1usQFP/i
Uo9sruCTR7H3eKOGDxP16xbe0QSzqvinbyRZk3ZLh6LQvkF4qYh/mU9KAsMLhjtg
5YcBLAHaq5ZeTcQ/WDH+oaAPJ41tniM+K257pSDd2txHCIi1S4HDrUQ7oAnThwrN
mb5rUygTlCrbHkwdorB2SMOx3A9tFJvwgy6dEms52KruhYmSsaPuPa514O/CKvEN
j5CG7WmtodjVQ9VaYOhYn6mj/NptLtkmUwi1kN/iUjvkJ51P/2UohbYOEN2xIo2w
9q9lQnjLicrrJwVxwggEtHYFGyuXkRRLNTe985CdYmFx84YfqdccSIHHnoBL0gTA
Aps5PHBLSMu0IjZGnvFz0WcLckuSSwmmSeZEMAEJTXW1QbqIaqYI7Y0idb4Qzehj
1E47x2/iHoHcrYb0Ozt0y3FmxUwORSABnzwKubWhXJs0NvINx2bckKwrMuVGx9PQ
4buI5lgvwvFb0xZKOUCDJttKPFRENd9WRqFfl6S7Vo4BwB3+nyweEJ0u1Paw+YkL
l0bedIP5bXH/OPXlmclu/MAGdr0D1AvVbbcO6enkRlRKDvbRvYZHuuoTEKvI7e1B
h2OBDLDzVAuz7gwnJe2Bt8yrNVl59HjLb+e17dvabHEQ6oq7tG9mPfHSs3GYqXHC
F3ZGVCnQd5qONI8gO9fZ9NcnWkjGqMG5zW/aKkoivFc9JQ5GPSyVhSkmFng+DrLM
nF2msA5CcfVmXHhVMJjAnAnuiSEeoq+eXkrnaRu7pjFrl9mhfrLOfxH5N3PtSVFV
U7/W/b1FpnNhGiqWZApqUgv47A8rsfcthcuFpqdqnd9RRE960fTYSGmLUoCO7ZpN
T4sJPJunQbv7mUSAEA6M/4fFEgGXS8dp5R5M8TIlvfqxuTqP4KV5ERm+bve8WjCo
Xyr46k/AqkhsFH4bsfrHxj3iRtcuV4sTc0D/D+D/uI5T6HgAzqNhaTjt6tViXDVC
FtBDarveRcjwp5TTIrWNCiFKRsLzO9+qnWx9PDLzpCqCTvfynWl54unSbeTjBR9U
dt/fn820bnk/6UOEaVuJIgD/bd2jRZyF/peCcMUiJyzWRnU57Z2dMRifBPM5BVi4
dsRR1YC37I+auhSrCFdJS5XSch9jnrU4aPMFNxWPzDT9cyAw6z7mKiraL8018HI5
Fo7qRT6q0eKBA6hpnumTjYGgzUXdNmL/ocu4TO+dOiHedfM6De5G4n5SaCsUjUsv
Ax9kM3czc3wf+DIoaHdjLNdir2dwW7LHAVMCFwQ+FR2GCmhLvargvnwZClaFRxcV
CE3NpUn6KOEzz3bv5D3WIG3qogCckB7BujwdL3f6SHGykQbK9LdG3Mte7qyxOv0m
PbKe5rmV8adZ7N7iZvuqbtvgn+wFdkV+wrwBKHuQC6cExH3X5bInFgF9t2qRPQLx
IQ4lOU0jNKD+8O/rxuq3NWN4RIcfW92KtDDKSbTBbU1GjpdQ95IdNtL5RmNQl6lA
pIxXEjf7WM7yETEXYxpWJbLMzNlKjQjRMysmlWKDdQ6hdF6RM9p92Q+91kgV5it3
8r9JMX0U7oP7cEZPOuNoyjumQLGO5jGcr0RTT15xTx0xF3f5sKdQ2ZshOtoSkHk1
HSP/pvCHWvy2mL8+b8lXgxLXCL4wbYIVfw+7LSt011JTBeF00nLI7lZbHlPF2jjC
HtHJFQIHhcha/Q08Ovj+FLbOyi4drdUfVQzLUPZ02tVMuT+ZrM/aXMhJCk2fBkc2
ZAlU+TvE5ik40kUb2E+s4EQYAwTGsDFNAtQev+HnJoV7X2KORRSMs3ILcoRDP0ub
B4S4xmJOwzuQ62Iz49o6M0hRPE0eUcp7mc33iNhW5MObEdDBJhFQGSc8v28Z/OQU
ofMGYvw2SUmqrFbLghfru6agffrs5A1ZiaaxF6SypLP3stkGdKfWtyONrOVToXML
fX4E610g2/rogU6h/fkpzUwu8ZThAa+Igj0tKmDjK1ZDKKGfZnlr4UeSLcK/VcSL
7w7q7uMc0ZspvJnPtgni8O+3su3DTIMACdbE27KaSI15CZ8dmjYr3uX/PKEBfwDI
gFCgSfTI6L/2FvV5Rz0cATEhjq8VD9mttyUQ2NvM8gbUDsoymcyQ7FAgfBqkR0rr
Ds3vKJEkRL1Ady4JEMQO1DEtDFzxEI7kOUnCGI5v02bqha48mn74ABJxT53tM506
sOal3cyiy+WGlMVFJhkZtYOEnVR6uDZ/X3KuHJDWiiuhuMlJZ74VsOKjNm8veGdB
wKlYsCmwEm9j9Y2ORs600XAoYBaQDHQ7UtEvt1hihcnwwThACAyV7Kr0gz+m+Sbp
e4LYUjMEiZtEQil7N08YyXaaPadG07PfK/t+80inut+Km/SKRuloqvpKqmu1nMif
jtyAF9/A+IhXWC8njUvewvPbSQJi0HOUkFUinzcC5UcC529Df8+FCBxhUqK4+8FJ
i7nEskFXJqQfi9tI0hJfICrPhVQpfwLS/Hwc+FHGft3EpAOR1xx0Piq+1AbWqoNc
eUM7Eh15GB/DgiwZi8QmIoErh7xwVT8RV5ulHWXh6IcZQ25GABIVFqsYhJlDRy2h
VeYHq1FKBhTuAmFfrG3IJUxpnQllWnWpeR33E3J35y15IsDJPlV37hbjxtBKvYff
/pFLU49HxlKth8M33tKO6BidFF99K/BdArxtm2bReOnVGGUW++CXAC75CkJo5T9o
xMfjbd3Z+pgouAM60qE71zFCXH4DPozmgh/oEbwNvPxleHalIf7/xmjJG0ia5Pr4
H99b+moegv+Uy0/d/j20bYEXXxfszjO4u9/gUL+WspvJi/Tlq/lyb7bEhPLtj0xc
Mc5iTLsfzg/AbTYyaE6k839DFDDbZtINwcaWykd0H5JZsmdx401nl0aIqSv0ANNR
FZC8Q+hYEKLG/rx2Kn+daj2by4cmMGhgZK28/jAvEjAc6235NdcBT+R0iMuW8pt7
L5bPpNU1PPRwQ361twKxbMG1o2FR7OXTaLyAocZt4WeID0CSgF2cDwg7tJs51idl
36FOLbVWuATayniXRH7q49OuNZJOBCs14oRTIjbrQl7xoNsa/OC2cpwNBHd7Sh68
zU4nmJxjDlO1W2Ivk3qBhiksK4mhROvqCXSVM/XWUw2bFYY2j+++gGViO9CqcdsP
FWrdt6Up4GCa/j6n2vRVGgvXLH2CRJwIW1mT9b4kYLSANTwJQnrNiHovA3m7oVsC
Ckr6nEQzT+uAWoRUfq+lH9pTcVbHkZntS3Vn6HyfaXPnyoJXJwjhGpwe/ZcsaOmE
4ebHTv2e4uiTm5pFCLsRSWjPBHFUZq5CvpfyVf7IRBoxPHlfXDkQ2hP8+Roi2fK6
7PI7ZagLBLSbmL6OAi3GSdM5CUdtKsQv/lJmYemOYfru5NWviNoJJYf0bvq2eMyR
u8ob4zGtU3Fcw/X6tpVp+dqLBAqkiKtyFCNnImjraYQupa5XWom7nXncx4Lbe4hR
ckejH0nh5dpgpZW7BW+EsRNbGtEJFvV6rnMy5xL/ZagJrPMEGBMjtfJUxroHtwc/
fI3iNpU5cJW818VElqDN+vKlbUWJvFJdAeLqjb58c+HkXGMLUgCk/F6vsEKJyUdd
Si4TnDu4fFq9p3/2/2JhCTCwv35jd9xoDvP5Xczd8hkIwfsKXFnSxWxRbB1as/kC
5Lai+qOGeQ/jP3ZaEc9177wgx4M9+hsf5367c2sUqPivO74coKIWv7Jvb/Fl79W/
de/h/zxLI9Iiv1aZkTJuMYdad3Ld6t/wz243h4M83j/Vs3E/ZO0+/rt1DOZkACqP
OqcEv145e9mvdutL/3Odi0TZZZNP0mo+dmSmnolp6I8dtGNuFub+trKCsAf6HINq
FG+4G2xLY2y6mCUbw3SpFRivhjcUjixNC5C9o7t4lBW6vtmbpjmc/xzLbE8MWvKE
RJRRApONOhp0fUnBRr9SUjdpNsOfl9ciREHy3hqq3A9y/F71uw6CpiRhMiG2YCpM
86CT29zTfJaUhrYCt/8rh8VBXZQHjX8nFXyx8Y79mPc2eGnjC3nP4CFg3jhcILWb
MoeMa9rIqkfmukuU+6cZrl+NgXHAj8bcajUHD19zrGI0qJJk09dDxKz2p+jr5AQF
Rp/kM8jo0tEaE4J4uYm+UZlQ0tM+9lznNWnZj7deMZquBCjMjsoFmbEZp7GkVv9w
vcbyvMa/zw6mVEufIdV8YkY0+BQ9WbkEo0BT2mvIKKHOTJwIDB5QbmdH4YzxUVZ3
YiuC9T9IEMcZeng6pXYps48uE4WGoyywtjsij49otjOnWx3NR3MWQJytb0N6b0+v
Ob046pblKl+Q7E7qvPGVsP8od10LarSOnBOJZCSJqykYM/RhDsl5CPGDyWoGYF78
k9ru/mL00ve0a9FfWcFTs+HFk6DB24NEJFa4mlOhD1W9POTNs0QYTK9H11tEOuJa
OwQNwsGiWJEHf9wckeJ0+0eELpXUsifYncYKC6yzNRSqmUYBnzHbnyu/dTybMhLk
KO/mBw06tdOIxG7T+yxzjjw8rYQt4LjibHKWO1dpCByNzCITiwzuAXxRSTg5HypL
xcPdVoECumR4Q7w9cYceqqhQw/j6YHJ9bKx2rC6h3ohZXfyfSAe2QJ7h7YQZcsjo
rxysumMEK57YSEoxPjOk+zbD/MdCzxluXnHU+fTaIl5PF1YrYGWNpOHX44m3rbwK
sicNMRxcfmDesUes5MPXXECLNabPnNxCt8MUerwECD3wk1p+TQgzaph3JXJb6JaY
LC/Z5+jnniB8P/7bc6TwaAnCvRaI5Vg5Ywd6RlTdXzLQ5oUT9c+5xFbBuTxbuGj0
MbHI3QQMdQdT8B/x82ZebFpyz3Wgo1hVM7EK9yhJpiNNz9HH71Vm17WJn+LSvAGR
276PRFvg3F4E0G6D8hRc7rMvL7yJJOWm+yYyWYGwAOt6GUS96EPPudWUR6dnEcCc
ePi8hmydXuTmZbjosf1lzVNDzkD+sbjeVRRJN9F8NR7G+pO81ZgjwtY6Jdf/NA9q
m5aThLWJa3YBbxfVCk3+pLylq0RDm05r11lRF4UT2O960ZH2NuI8hiFK+vuOvEqL
XMhDK0GEGOrjVwrw3G6M8fAQUh7zEhim5HwHa/ckhEcf4tQTbY7lIOStLiaXyVi+
uxDMmXpu6cMPV2z69fCwJbOlkUpzEJ7ZhILj8IcDaCp1TjaFSw4hVv3i8HgzicVc
oV7bRnUHea9KO65liP+R5bDoRRU0v1n2jgmy+eZ1H9RibEtk31NDnw76VX7pfw3f
aw+3OU/0sEDAU34MbovvmlSOczDyLd0qA3zj1+ssXTrICnJEByQk4hZH2cvxkbUT
hlZ+MaB4Zcx9SvhpkxukmO2GKVOujrYAx+31e3E5kaWBK+iQiCtv4vtT7CGBFSuF
oZiaPoqG1HrauNrNCioYoDTp6ZG+fTIwHJshHH1Jbynh7RmIzPQqe3HStgSU5lMM
smVePxTL3yru3wrQPQQy7EJeUkyDVox3khdqt/9Hu6r5gG7WAbM6iThBLGStpqLo
qzmss9hu/nXv9y0/jEkq2wazSv33FdkM9Fz7d4KtjWFAET0vJGIOm9dbK9r33wtV
XhWRAXirvseCEWwaoRc68KkUemvFmMykZUhmOKffhwjT69+jkbtOeCjUzxtBUXWz
2rOQ59/S90sTTCFEJgPOncPFzedoiaC114N2sOxSieOQ5qWfah6WA7Wj0EWwNzzv
xp6stems38ZP9k2d6Cvs1By5dHpcPGZvlXKMi4B3kS7fFUd9ELOOUGXG5aC/f5Ki
53y40spB+ROvmomXczamzo1kq6PrMWHaZSmj7jemrIAvoNsrKeZIy3Mw47/jc+Qm
mRbVMGqzfyLcsA9sYQ0Mh8j05IuJZQ+AfRlNEQTSCj+BdnlkSEuYb9lZdihaDlrW
hYfhiU+i5CnHvlfLKsWoxok1zGLhgxiG2gzd1g8PnjTIvn+XOvHYCjg68V+7EKvP
vhrmyhCR85VOyGyItpLfgPc4WRPZBclTVlf1x/F7kMETuBf0uHxg/+n2Nq3vFwK0
MSmAT3Rd/4pphjqOzu3MT6MaVcJhyzB6vRCtFIQsEDQ5KuofiThsnj1afv6HWi8v
dwSrQYMNH1wgMwcq12AIoTgJPcElS91VvFbGbLSnUgNzedr/zzr5w/Bo7TcgJWBv
e5LJQ31fH4c3jFBc/vLQr7s74yF+HDOaTuOJDcbtCJtYsISPr+sVgjg7u7Hrh27s
z6yU8/QGH6eusuzkC91L5l0xyqJQoJhCsa27z/bpBLo69Y/DyADrsQOPIPymXj+r
+SUJQn0yM1/NXTAkdFbIwSNuQI9Ew+Rle9j9aGa/59V33nlp5Rl1ifip32fPNXow
dvWZkVZLW0bV5+orQCPSwlkBBGL6Y8lCHdOqdFsRn+DoZf33YDIDioMxZ8WmcNok
jSUYon5IHdL40xGwI8JjjbeSsQ8SCP5ki1lTWiqXZsWWwTeYUpBwivl1aglW0cV8
oiOgWCyILEe4nJXJTMCVGO0MGG2cLkvkyP5CeIwIbl//nk3fFS9P2ZJ9fHGChdt3
mW8vFP5nZwR4Hheli9OAo687R54Djhwwp7FCkA7Cr06qE8Jwm9mdmM9j3i0ut3ui
6pBwtfeGFZ4286FQvHkRO4LQFkukPTcc3Rw6uuZRDMuNWZeqMRed71eW3x/idJyb
0rmQsv+/436Dyaaz67WHss/Wm+jPP/DleQxW1wem8z6tPrs2snIoTzAz5iWcZIiB
kdzR4oOWqu5ZO/TsvGXWsrUZHE056sLw4VN9R7Aa7CN4c+aY5/F45cghJ6s2AVJf
YamMDtzW24QKa94txfngjzCb0w9DG12r/F2vqzI6cTwY/9ODI/uMYKR5krnYZOc5
TkoZjVpdBwbFXqbYgK4VzgeghMDMb/FH43sJ4Bn3JJ8BTa58heN1L8axAmtiynUH
uHh7soEZERb2fAuAA3EFwFT+tY+GtvB01GUTE/jiPFKbB8iazxB16EE3WDXG0pfn
ztPJeMMyQMb+iNQfXKGSragv5VzEdJ4DEgncUJ48Ha3CDT6YUyzBFtFi0BeBScHm
3Gig1TAOox7otuEDwDda8gYpuHb0WfxRksUu620SIAvqWaWbZ23Hs/9dNEV+S/Kd
o3R7a1JrJuvxbzsTv810vU3OitullbXoFERxInCaeafy0xYd2RkNptH+g+mYu8hh
jZ2GLJNc2ZBE73FcBt193hirRufRy46w4EivKm5ROm0QLXzj6gZBbt9Ht/4zBp6d
UlbxWR9ADdYsy7dIZrG7/4xcqXzmk6P9xs/a1spt6GJpEPgf6a7viAXs7wbO/gC6
ysSuR5O+y1IHmiaeW6LCOghayLLkfmnUzZ0Sy01NIRaRZRLd/nnb8+sQRPXF9nEP
sJmdFoOy3NDXNh9vwKSoAaXyVjrKpvKOCk61Own4YYts8QZ0mBN2CgezsJm7wbcs
itKWurEQ5ilhLH3guoIcgWYfhESQdO2P1ylS3tKmrmhzJ85YLOtihUyDDq2ptO/T
TC02ArVYLl5GzCHJBz7pZdBOwyGbohHdeI+oWhVhQPXfS/GdwVvZVNHvak4+1yiw
dnNvJbNE6BkJehPgTe936av2U2Xt6eCIunE7hCYUd/tQ/SJ4udxPDsSdTBW9IX1y
eEIu6GlXbkkScupKdm+d1t7k9Og7934vCziu5AUKAovLsk5yKTd8Fws6aPXYjZSv
d+RauudjHpCi1dTnzFknIbPg1/a1ORyGj6Jogg70T0d/bqQgq03YozItpNAb3yA0
QmzdgCp53esNxcctQEOyL3/y+8Q8hMqdel+6E4pwmFrqJu/Z/1I8R7WuBwmiDHGL
OdGd224uyKLjBZ4WfZw9l+ECOdVYudzxAn6tceSpbJmDCgCjumOGL7G9MsoEInu5
G8nMMll9pEy20triIFV9w85zjNNXdjG43Fm5Blf91hQQ6s+lTF0t8hYEG0T7wW/e
GzVDDUT/n5CITeL7mmCU9eiqFItyqUxq/YPLnnBIc/8ID98iDV/soNj5bzS+185Q
4rjFR6Aa1ZYFEfA1i01MPP+szGJ//ESRJuVKb4B6+133SAnSMiCjS+K9JzF9+5Gs
tHkyk9aD9wMqhocYI5KXnrr7rOU8FVXaf1tHJqNUgcix84+kQed1nbjsPZozICrW
BmODWcPIN/mgyc9hdsFPiTJ7UB/rfk6m1xxC33xU7ZyP/bTDFU3LaleUJHeEqyiy
j+75z7s+QJSbYJUaZDOYKz56AEEx8BO7kP9lyUcC2SjJqdDjybqs4bBIobCv1/sS
QimFm6IS4q34HsZLl9ct79C++sxSK6VEvLrS8m7pv15lSqMJRYYkCSJOMwthfIdS
LVNLaQz8h/YFxRNpEQwUd7be469oYo1Jdum6531CbincznsnJT+SY/XnA9kNIr9d
XI9uC0+pcpftuR7ZkcMXhP1m14xG4gLwOib2N3OD7pGROgnHqnlGI0JaJPjUeJCc
LyelRg2Nf2QTjcj1yjI00U0n9SrmGYMpKCIiuEN2hiwB+FQWUpojtjr+qDaRr1kd
wlemjWZal+c/K5QzrdDxT0cs0G1U/khZrvG3me5pp9mRFX6f2ynwe+KbwBR+7iYg
Ki1v1Qw/sXGAMvIwK3YAHE1SJSQNlG3oeIVIVJqEC4xSIXfsY0Aq8fzCfuPAX5DC
unA4wmTwCp8hzfdNmizNlq8N1hK6pBLxKzwiPQA3Ta1Mk+qhwWNurLp/2fw1d/Xm
o7poLXLobC0U06IcgTH8APCc4QBWUPk7/QJeN/QVsrIxcdDEHlaeBFzANuANV/+M
0m5hC/JToEAtSyC0Yq6NPC0H+vy3ID6r13fleJQfmyYkzJy6nUOEWw4ITHZr8M27
LIONJnqqNqB0amQr/YczEN82hoSoJnwyQ2+in59r6BJRI20s3K7CLv4yyYT4QsgM
BePf1y9Y0priU1wncvBWecGq73kcpywwhZ6nQa2yXMz6x3ZhXiD3QcvFvKl1QPSN
04WGoPE+Bx0HVkWZvCtuMiCTililhbTuxEy8nFY83BE9VEFsWlhwCSvLLENFTQEv
bjI0PKRLFqj2qhGin4Jm3AHCy+49AnekepePD4ht0o4ox+kk1Lq64QtxpRDk/Xz2
OT2us4S3P3UkUwquP8vX0YQhPy/d+9PVP1BuJjc87WSsXXfU9g61TgGssGgnoZKu
OtnMJ0BOo6gV+xKBALl02P3liurccqUrnT5Cr7r/DI0rqyD2EH0vNTKwjPU70CQP
k8wVTC2+9jomjwWnlZT/rhe9yk/aTde6/LvWNOswHEo2chceRk6xuc6hldYp2pa0
4h6Yg2nIr0FFHJz4l6ntPl5By9XrxK7w59jXYu/AiQdtAHvktnr8gIqcBlHtR/Dh
ZhDwdxu/V4ZrgI7YBmzrDJityAdFAFuxPytfPV/UdwYmkSA/60HqGjZpe4DL7bz0
ztnNHxO6ZoUX/8CzFB+OL3FRZpwYJnrhRVTYr9Gupi0Rb8mkzI/2IrI/dl55oGWz
D8T7vfvJsUeX0aGaXA+tIbJoQUtQROGun9BO9BE9Pj+5iP7TckmO5WVSDnZXasYL
gpHVMOXv01Ej11XGymnPUXllkBaU5GR6lNFzHIuvetmq3fnsTIv+SP0CRHep/NJu
aaEjj8nSy4yOTWyNY/4IAXC2//BSRVTm0iOEQzSbHCkbVrn/ec/+foZ+igAJ/ykM
Im5d+XCkHyTPOCDDtOqNzFfKjvXgg53IjGl3Z99C7RlxKgzbdJgjgQNR3qnHYqMi
YS4MC5YMbbasrLIHa4PoGE7GQi7389Ax8200FLyvebqTxajzm4+Awm7YwiGy1Ylm
uk1tNyHYE+JG9iw8lw/kBIzDCUwxe9loRPoFwxKIGsTLqYYQC4d2fNJGMlc0bEKC
BEK8PUffujq7QsJa5LDKPFqoW6f/LmyzitbV1FcE/AP+t9Lya/KmRcX4gnj9kZ+c
yMqmMNdXZfhaW7ae3lP3O/MxEhTApUi7z7+qXLx474nfShcoJpEngDT/HC9GJ5vr
roBfLOZyinUmS/gYLZJj+Cl9whZvH1i+vevRM4QzKCcWfy+En+g4tUlJxxcn3iq6
Ez57xziP3W3gYU9eU4oQaHV/MpZwR0hjCLI+N+rpjoj8oi6+OKH3mgFtxsag0A5R
VjflmytJrTGZckhJ3pzsk5ahq+n/B0IlRyZ13vgzSM3NICgQ8dRmoQF1IoIWJOaa
wHps8h76vnAWNss/Ktx4EJUNtcf14dkwU4EZal4fFEdzDZ5F3YpwcIvxxonmAxKG
f4rhnnBEqNZ9Swc+4elbVCjbWMSwtNfIz7tNNpTFt4WDH+6BRmZH99K2kXiQPNmX
OihbEt6Gism41zpzxVYCwMUUBATUlDZMz2HSsR7XLRVEsgEEUq4iTq53eo/q71UY
96SQwSSq8CJes5/Le8T1atf9oO1Zi4ogPvaVq1qSrI2Ew1Smwl5VYjQ8Gs91t306
xMh63ax6mJiH+s2H+2cehoOaYcpU+MM4PXLdAe4TUHHhEUgh4cxckov9vgKzAnqs
DtyMGLtw8qDSRwtS4fjmb0oNK7L+fC1/S+skk9FZ36vJWaul3++xyID9UjbowdbD
LokEQ9ek475Rxtr9YNLCiycHkquX+q+JIWqG7v01h/wvTOlVO2sitmL1qpf2kg2S
/R0y+zzzA/ED1xZWaQX9FTNhZFRxlFDvvclkWGaWKyDL4/8PgVOn5P7PCCiplsBy
9swy4mxhx9+zJXUdMRalQHJqkj+1jz6cGXaDXkDFToJs+GFD1zewe7f9Yn5awx9x
zlzsfkKATFdKA0HuUAQ7joiklWoWw1wHlu/lm3MJFnES/BswpoRusa6Fb7ubkAKQ
SIfG4VL5R/1X66Y3cnMyWM6zpZrzwk0Et8p0HL+f2HYuEaKwAFaYchxz+5pojPHC
Gj1Jv/M4XXtvnuDBeBMPwWudxP4uMUOLYdaSvLRfcQ2B9M918e1cFH+2EPa35I56
AnFwc8x7RS25b8TVOf9FgZX2SyuD/qy3Bo0DcVJkDlIDxVCsAxqGcAU7lih8SpHk
IoN2kKCduns3n36wpH/FbyOo/CLpoAQ1Ka5vIbgHwFbhxbA2qTadgeqTYVr1/EDE
PuHZOtDF7jLbWDhhJ/3w474lrixsgpP7b4CA5yIjHwfbLkiJeZOZp8ONAipDFY71
yRLm0TkXMN954IBVH+scjvZWSu4b286xaQ9PPgVBMTCdpZ3oLaUFvJR/Nl7+3t1J
mhIx66wC86MOm+fXbURQ1bYlXBZfvow1dVHZZ6wqPVt+Xtm1CbZGao/DNJH2T20u
b7eDwQEvQSJI8X4v5avd+tL3odiKze2qnWjliux832XRvBfgQDR2ZJRS+a7r4eZL
fT1dKHqORlv1YovWJQCvXrfUDIhwSUp6fGf61rSS/1s+Shp7ZwyxRpR+N+T6mxsF
RGRAx4O/VbWL7vYGluVD03Rx36H8FMZAJzZfAdyDr7QnhAXBK37VjgwTlsRVdkwH
onCuF5Jar5etqPv6KLdeXtZqhe6d8TSePgFgQ/jEbw/lrfT4L303iFL+XfBevgaa
QFqWqDGE9bQYkdjsnryoQ3v0TCVrwSIVxDY/TYrJOEHorWeODiRUhk/6EjuqygdU
8ziQ6Kfx0q+4efTRilOv7t90ct+jU+CELocZxt3vCamitSmgtRmV0YfeQcxY+uDa
QWt116OTLFJr3vh5RJ/EVKV/0kH2HuBYkpGMn2IYw2Uqjs7zvU20r/0CbP1HdCju
qkntrX/WfeOPmx0Od8L3bvvXyU0OukbgHej5qZJgbakIBKe3p4hWyDCjQTueWJE2
KVDVe4dPpuCKOQ/eNbbjcmIfzpO5cnD7cZCnTuNEzDTAjz4VrnWFAENApDtEf7cc
U6yyckaTeDgyol5eJG+27CutRHyz7QhwIhrwcDgQhRjw6uV2hsWnjoXYrl354n/D
R4VWQezTr7FrR916uFr8LUvuOtzThd3Dy5+/BXwKjded0sk3HMg++gxqhiprEOXt
4gAxjJTznHaGnc5PHEm4EgI8vyI1vEw6VVBQxNZ2KTNjPB3u1SLNLzc1HLBXCAz1
bv16hCRvAzbSKCUqa5nKEpmpLmXN8KOFc1eWmNmQHFpfc/+hrL7C9D69KrWDzr/B
Q6SnGW5AKnyJ3v7wkmOsNBitMn+nYOG60+ZxhOQJTx/9eYmpue3C9Mf5Db4hR1da
8fZzdd0uvd/GBdDwvv9Meqqv7F2tPWVTITl7hPm5SXEFEyjutLE9nIkr+UTM6ILZ
/vMXPQkIK//6IQnKGD3GwVlsbc8QzugFkawEShW+B3dRHlni2qMc7v+/cuDDKObH
F/te7zStABzhhkVSEAYJo8zYhpvw9RCQltf4eKDXOgFfo8rO80Qkb+xwlO3QuZmA
Hb8SdTMXkrA+Ds/+nVPx1KsisDBlcUakOtK2HTDrcNNYwdOaIZX8luClRL3WICPd
SouwIY2Puvig+g/jyvzwC6M3swTEiu6EdJ0lgrDANtfkq9zUgEJyCLHypGn01sKc
aO9s5k1UnbxITwdbtJ3W+r1RtffP9P6KyMDavpBC9XnwPGOd+VdYPIeZhTnndhLE
8wSdzzobdfEfwxOjd70pvHXLKYUOKk6nQsmInfs6JTKExrM/L+EkK4TWF1YONVot
N/aKTbpXfe6v+NEivJnl6gPyKjX9aVxtX9gbCCwEkjlqmO4jYDG3S/MdKHj9YfFl
L9F5wxSW8raZf42KBoXUgT5VaNTIdEXeJpPLDuaIvPXraRBvh3hj4Yu6/a9Lqr1x
LeUFuaqZhr9Ajl+FS1FCiCJYCv+2Vj8NH8wt/Cc5nnrtoGk4ga/M+5y74nDpPw7p
YpwfdeNwYAYdsT4Vkynl36j+TYupDClJYRHfSAoXUGHr8BbMhtSncU7bb+13lkNB
H6HTptJKcMwnhdcapAT0AqGyBPDwAKikVzw2oVEJ+5Uyuzbu7OxcxKcEkUWHNLyy
WzNIyy9pAcag1FbJMyyrL38X2aaMx1JvD7brBB8biaNEUf0tD78bsckuOpnDfeZN
OLxhwQ84Do+0ZzynMb21+3nQXjmyPWA+Lz/vG8Comraoob6T+/42PSknsbvcYcmv
Rx0NjFyPC9MJEKHfUDd/0Twh/KtXM8teraWLQBghiHT8wVK5b/xaVuLSide1IGVs
pznS4EMnxL4uJxWFhC8oEfmyGVQ4AZUczo3V5HF+Ndu5RfpI6Snmv+lyi358Ab1S
O2jfqfUZ8WxNlNT9XmvPDZ2XB+U01bdzbASIIobQC8KXKwCFzT6t5wfjLbDWneU6
twAwlRK6oxLw1pYQqyafy7CntWlDuqGg0cO3CW5hydh12ka8y897v7GIdB2MZqLy
ShH2f8f6hMV5aOKAii3CTov8UhEzbh2PTydhyUAwiPZTmyKiCongWmavA5vKjw/x
0Z4YX2rvf1vmZvUxy13g7A3dPnDPd+0VScM8O2p8Bn8hOdobgfTx2fn8uHM/8QLo
59aqh1jMo/jEdxhXiaHgKJCfzomOS2Hbf0RAimQMawy3npJO1m/d7M7aJJybmexk
FyyZMaw/836dZZs64skSYCNvaoVMZe2gFowzRtBptzWd3GFM2T2trw7wWD2ZX6dm
CR7zxPZe6z5wdUH3pDLokuEOJsPYUj4CnbFl48CZrJOmr+ESE2BOSzDgvjlyr3rc
Bi1EA3f7AJCZQjlOtb9rT02L8t9bqOF+gcIOu/aeuYg+Yw+uMXQGqqdbF+gpoYPE
Nbt9nEOMIY6Qj5EFivKqW66p/okLE8bVg9Vrtid6PjTkqPGzk7clnmeJPZ9ED1v3
i3r8kOiiRwZykeCWTniRL/1v1DtsRoa231tctj+Ueh8O0/59MPPY58TM6Vs0ZKDJ
6JcSiXRkHnsfdChJxTYQ7shrXDMYheGKsQwc3Y/APxT7gdUI0TY0A5EW7wXRHIb5
WI+2cHFAPSMbxK5piJsV1wx97xo7G9lU7KmkUfTa1V94HZ7LUekOUSkbAQJMUdkb
PDzICktoVPgpLYn+ouSlcNY3eFr/Loe529Geir6ABD26Tu/v9Bsu5d/+ggya4Xfz
XQ7WY9g++kWojghMRp4XnnI/A9A8tMwZeHiPGNv/qUZ3/8b2tEzgGzqaVMj0B281
4DWeqUj68qYFepqekoljwjMw2hJZ7bdZAw3pWxJ9vu07P2nppvUkjr17+RI0cp11
CtRsBPIgWpNjBe+PuozOYr0eyAXS+ZETRxYh4QIFpz2Cip1R0EoSJksLuWQBs0Fi
ljWYmBPoSeVhQp4DMPvRAWyfxBGq6MbckkFqUIwcPHJfxY2BL5GlGNE6HYwk/HY5
cK6gk5Qf3Pp8SPYVhoNI4Egils9s67Tux3NsMsaAamnx37dO8cogwMms4+9suCo+
QO4Qq3YHe8RBLe/eTRh76k2eRNRhmo4C+knvMUa3aDmMwBxha5kLnV79nqO34PZT
j0m3asOZyWuz6cn2n6Mat6Sg0P/emKtErXg95n0Sb7RfBX5ZPFvS2WWSV95Y+Iml
/tvbSC9gkuTlx8CXXGdsX4CQlFMEucftTxQ2dmyq0CZcHjpXjNF/1+yQukav3Hfn
j4Sd5xvqOb/tAk9xN+JacllGPaduTqxwKKNbmkA+DrLjZ2n69AhD2py8RBZ2mxfD
5vr52IHxjgnzJFp53YAiyzBWRBqyVNftkz4Y9k6f2U7Djg5eYVxBhVQXD+1/m+ys
DhzdGhIwJY/oI8EH00TWmcUKOq7hHxebNJvpzbtkoCt4Jk3T/JJwq1diA2NFpz05
Yk74S4bKbGM5pMl+zPubJpg9+abwZXuPQ2tNnTxOUN8I8yM344BaiMSUoB68MSpu
dzPmZ14HDuyVtyFKQ3EBi3r4yZgUfi2/k1kZkl8LFK9Sa1i04rIEKb7Yjhw8Z5dX
TlKPRB6D6ZG67dsBJHXoEznvP/dFeZrGdbxiKaTSvKmSKV8ZVLmioZmLSw8cBUPY
UDuAT2cNAa5ZgPCdTPOu1PDP2SkMTUGoHb4Dkdp2uSwjhHBmHSM8qspgVVenD4z6
JSnhmKtbNi+2XQtNC6nzJ+RjXrGjudFNnvdS0/cymHyIpWEUCHHEb8QW7yzgviSq
O0WYTPrczZu1zJdnCd8mOFcfXzCYa/xTrSx6Wdt+Z314D3mzVRBLGBVPy86XFb/T
/BqFA7F3zbYvXFj2wIC+163HUIE/tYlDvgAOmI0w3xFAuBWgMyunxxYx7wlaq5/j
Y4xE7ovAv4/XOdpo9CfusiEMiHZZx65yh4n2To/lsRqJw1q0HyR89qf9dUKFun9S
af9qAJSfvzB8zbGUr3eehSFXElcFJKtxrXTdG6zzvowkYZcpxSBSV+m1CaMurXM5
1mEKp9ANr/3V9LHC5E4SRcgejQWdJQOYqgbZHa9k75LKk08uLN0o+KQWkJFUC+Oc
i8rDG/kuXbU9gfaW4sozlZO2ucJKoPmswI/0guyA9rh55qmy2DYm6AbinwcWqJwY
yf605kO/YtcBPMRoBf5pdp4UKEgOlmAx7NMxg0XIYT2QAMHX8hfIS3hisOQBMO4G
Fp3443lBDcjpFzJmPcpNn9NphhXaO1tPBBH1duWiKcgnSbOyr2EaXbykuNix7Vaz
GFivVFANQKKZnHQcr4VNfhJ1RcqyYCarb8obq2wdKysNSU0twyAldzQFF+YHHBe/
aYPCfJYDecrPsFPPKWtGZNVNZRCsCh8xtMscW21A8A+Ic/T1Ysq2IcBeSV63OUps
fzhWSx6rJbhRna9oT9LiutJoXgqEx+AptLW5WxFb7E3t5onTwM+/1H9oyCCjrkSB
2QgwX4GAboonz8R+ypDDtDOrWco4OJjp2F1FNB7gw5/2FfJGeoFREH6jBD29GC9g
4pgqnoZuCd2BCK4jYaeziLOz1L2aAYHfK1alkRf+DhNxuS9j26m/UWhthFWeiTQH
5KaWaIsAQG0fVhjVnRXdJYozvUUOie2bKMlWsN617AIwCfA4x56q+rhgeZJ1me9Z
0Rvc1g7gmGcvlXYtUaMu4luBeEc6AyQMCL+vw4qQOlII5laAMsQyt4uDf/CGRzuP
ESzAHk6ZSZSw+/IUzdGmQCpvV2cRUJCCAV3wg7nHiBm26q9tztV1CxRF+cxgiuzF
h3oQOlmMOHticxvYJ1SpK7dV1h7Bp1K4HXfvRuPJ3m7gV3rHuNNTYdn69zk3Q1Hp
IFJNhC+78um72KBQYzAeipnYP39Hm6EGAjC2DXW6G6SxtZSiAcU/olsEmnMQKuqe
ZfJnusFSGI+opxVYf//ndGhTNbJDrJn8arg9nBdghYH61iZxrK4UZ4WeGn+55jYY
egKSf+1Gcnug0SI32EF7G/Z/BpfqdYZXinM2/79BJ9rEVe88z8fkqP+I3c5PSM1j
8HWO1/cJPuOrb4BIcujJCzd04FU5bK4vQkLVQt9iaLemLRVpZWQypXMyv7mmBIfe
EpUP4FccAPA0jCgesIDSbnIqZ5xcHmiGxWnG0PyaXcPyqFGjo7xbV5X7J+kJCHZr
5C3DHivh+OF7jHUABLKrzb8NT9F2BMuRpbm2Q7HEYx2nJ3M8NxWHANicv0FgqX55
Psc1W5vVDtf0mzVZj456t2OAXB6+fGttnhJyKavZyKyUBUuBVbaU7nwA4V7yXriM
VBqHfxJ9Akzt+EYOfSnqTAHbw3b249vC+yhJTwuhglhSWSgLBAqJjcKJjPH1VTIA
H7qLZS+iVZhDff3Ak5kLVoQd3e5H4hbFH+E6AAK0PmrnNQCFzwC+/0W1GCbcib1r
jWBq+4om1X8NzHB6Yg+THdAVJfSDQlkSQTae2OTYjcF1jSlBcs8DytOStjGqSGvM
Tnl1qV3+rKPnGT7f72/xdfUuY5FfeyFyrFqALRkrTxE6RnjvHOunqpnKyvmS7eeY
8Wv1QI6EQJZ2MOE6FBugAkLqX50n+n3b7EDUDGgumXrAAfh/dFhxCf0c/VocGmjC
sfphpfs403E/habAuEPRYVgXWOaD7sbGSRF3geBDroDSrJQ6lIhjqaje2BKAezRw
2FB1bIM2t2nxpvAo/SWyKuvjIfWQ1dxfXpz1RyKnJc9PQRjk3UfK/sZOYzuIgi1/
QtIbHHAB23Dn/wAtg2bUF3lvrQYQ+gGHoiwiRZDrIXWPLugZXwn70phoigze0gHe
Rg3dV9Vcj/nhUWR7f90OMRwSjwYnYXDGyuzhm1Jaf9jCd2fm1hOe8rqdNiaHwp9m
YPWMmGCqSseB50QxpGd7bqesU10u7K8sPDPdqa+DjulfcJ6M9T3F50EPw1LnjxMO
aUyhPUrGGgXF+LSeEsTlUYiyc+bdoN2rricI+OhU/DOfmXlolxlRTb3HseY+TW9G
ksq7aS6Q89YjJHn1Mx5a0ZPY5/SP8E3culHrhvwtSVdh+TPTfQ/R8rk17yzABxlz
2j9DGQTbr6EAmhBvQdZ3gc9rmGb2Lp6CqQZGdcqNGZbqk93RU869nwdBm+ieL/AZ
Wxy4cR/6WhMfI/IPCjPb8UgUu8ldmKxIj7sJIyuYTF2Qr51OJhd21W4tLEIAQnNG
o9Irc9MPvdLhq/KZ93N62Fq1xe9tLLl5uX+A2o/S5cu1oHSx4xUNLPkpwFMjGuen
gnpb66x4nWCTCNspydOWeJBqEoWviZEFktHOOrMGiavt1S1PXxPj0SdJdSork5rn
K9zMDrHpO7d8UNdO6zZNM/81YkWxuC6H0p3fMUrvJiDk0kkUAO9p/M/PH9/xJK4P
NwpoSE2YgIkcEGS+dYch1vosYaanhyQV2KqsYBGKXWUHr1LAAj+9xpWW2zUMqigZ
1yiFpKn7Guc3G+MyZe1KLi8resG301Q5qM5hDvz2cyKiw0t1qMi/5AWEJ4ti82Zv
I+bf1ofh0j0DxrUgNSyyY8mfd82Ftrk+L/LqLCUZR/Oa99Gy+s3Hf4MB3iSKmWA8
piZPKYSTu0Taj4//DxfnwV/y7jWqL8GlveL+JpkWXa37q8nEp6cW6tsfD6E6Vp1F
NFm0axn0ooQZiV93qZH24T+yIQXbZNfYpSKby0isJfdjKi+RO78zXi6Vr/3VXm+y
2Y2MbYHd7OInuyUoPL8Pu9YkFtkVP9z+XZ4jOijV4T6u5RKw8ACRIHEnUI335akD
qYGX/HsF8QDqUsfxtF6h5IpIFoutamyzHWtR4jthc6BFgfFdfJMmYXZSLktum4sq
BA6ypUE81D2Q5Pkx7AY1vs+/hacCQWRINpD2sGGnIB5c79GcH8R3QechtI8zDdLN
8/l5z+Y+uvI2wDrEgl17FpLXQFW7+3km2k50m3tWj1vjTuPe3XxmV/F4I4ofxI66
P8vv8xVs60AnGTv4XVukLu9ka214PV7nYpCWS6paopqjufODvzpHIp6A7qAG1m+b
UkR/GzkpWlIQP8r0ggLmlemMb/ku4YGUsL/wVsMKDL/xFwN2KBCrni3vLc52XoPH
4Ydx8OmHZdVFlFKQSa6NJRQyUQVz0X65yd+cpX+ajaaKy2vu0N7+fI21J7Q/Q6Vo
HwncWSGUmOaHoELXMDzZfVlXlKy/139eqxXfTY0oPKUyP3Dpu8B6zVnsB0Z4vnas
/hZsRrkmwX9pentSAzqFi0lHXC5OJvrvTgEDt1H7sd3oKyRG+VYR85X/61LM4Klv
ars/d3Wnfh9uY7P9n3c7cB+TCSvvhr5ef4dGDSKaBkyzr+og+QXEyYctMjN/isTS
bbKPK4Ze/kKJVIlwJZtt/sgFGBNQVl56qB/0CMfoJiQTkf/6WLcsh/D5xZKX61ke
FS0xA1FcwwPNzVnwYrXU3j/lP11EieBVDCL3yagRtmlEEX2otc7jXi6CZQ3y+yMb
uuvlSLIRGgmckRGpAFDj+YBrY1To6g6x+GpqOgIRp3M1fuUAou8Fa+oUXUBjT5mo
2iaIATsoo+Aoqpqt+h7c+ZUmZktDEETY0cxqGdqcArxa85E6g8nA0DyHDCGkdKC4
V5h0RfNAEaIPZJWBzi5Ug4T+BTorKMruNL5EM8IUVXXAg9QqqmlqYra+SZ74bICO
JGp7umVrUSG3eTcmxPsHH0Chd6Jvvzs9Ed7p1NsfyhR6Ew+OvpTS2crOmoKxXpdf
KRTPOD9o6F20BziKsN5ggurmFkcwQA5GGr/uPQp/ywlxXAzUPUIl28sJ6OGH9wOG
nKOtCjTtFs0wcopRNaoL1dRm2agL+Zl1OyS/ySOna+Lbg3XXVywbhyGusumyun57
jSe6FeEHcuLKKSfn0eQzbmqRnKrFGnF0KfW8cy2WpEYnDvWmxb/LACM5MVKwqOrT
7l+bgMPq6QbPTiBL0DSTJAho7BCO2WD1Hp9P0ghDZCqWmYZIDeODs5bCg5FrxikJ
snKKYRBidRII1lL22FtoQh5CVt4myExaJ3gEHBh7noqcaX61srF1LVLhmydKkMj1
eO46zL6NYesZcGleRCWrvgrCFvpQv+j78BigHiAw2ktKx8pgZrQDX3hgU9YnsT43
HmByLfyW+fJoOlzkxmI22GLWGDrrQXuXat4Lb3jqfxV+3VLHJkdFl/IjklDSLVjW
PDmD2TQHPMeEjemReLW46D3GDEF5zSxcCrpiIQSzm3PIAckZGDMN92Q7fBhgwINj
quhp6wZErgNnBzYM7fROYjcGroxMbxosFIFqvVJzWqT6QX/4+2PfK0Dh6nQBr5kA
J0mM87hscFUR7zflRaW8A4f5oU1QIIE2DcD5VHuVAQFh+2OGRS+XkQvOOKrG7ftD
6kMVht36GrEDkwsaSFT27mc+rOZbT+ZP1/QiBD3T7cCcz7ygrMOwlt5vHi/8bU4/
QY+UxSUi6ioc37SQMbjAwxjOt6uMiEzQJ7pYXS0Ft/OU68RCjCD5Mvy8wgg58U3y
ItPfJvBP/1lftsMKlKBG489LGZYp1W3V3oSZrLwwXZUKblVddC5ikHFiksJgmgHO
339MmgXDckoMmFwjZtYDQgDfdV5SiLyW5ISP7t9pvvU2iJAGwNgF9fwks8Hq0xRc
qZc+hF3ilPoXB6ZNpYl2rv6Jpod0kRMy6H0M7q+1ni4TrP9ok0bU1MDfmNFXlPxq
lH7Dz3WrWYFK9iwynmXYab9HgyS1Nc9hgcVEAkuABxNXoItTuIF+YpQkwvmZrtXH
5xvq2uNCUXvGBFz8J172D5R+ZtJxTEP7msNdvM/QLNoLSQA8BkFKPvyoPvrvF4TI
rPXGAnz1V7aU6NBV9yyq6Twajp7Z+G5MvOEn1J3SKEcjyjJAnlVa8aNezFXCilk/
mbYo0OYgPhSyQ9zBD5W2jWFjZhJqZ0KPfvjvynThZxkTOsCYHdTg3HGBZ1LI33DW
NYgqmxFOp1yww6yL3sJvDS5GP70SADLvXSiy0mRu4k5GbpupMGTr6sSzM+IqGzXV
TzxcrHErU7oIZIId7n00ySZPvpRuhMFi+9c7PYyh0+uAy408rWa+hb4Z/gH8d/9Z
J4i2SJQRRtwlL7y+7sMiP0iNTUSJ8WjBnpiUk+t/lzMlUNJ8va08yJpX4HpWsZgB
ax9QjFp0+216j7MLWjnixxhfge2u/5VAW7jPWtRBj4+q75ZT5knS38AbQ1xAW8MF
jLKFjSIoL7LP+JTvcUi8LR+w5lrWtQ5IGRcWSfyHj2Umhrn0wrjG3OE/JQEe3tHq
9wK0v3vMkv6onpujE24TR19UB/Efl5848XZC4R9FLDmup1jUfdMECSSicvHGMjI6
iDGAp1EO6MnSFbHP5ae2aX4F+mReEGHZ6W1d7dnB17OsQ1IHLK67c8neE/XBAGjP
Uuv7kOFQjpX85iFYwGSQCljAlD3GiWITDTVWkwf3Wt0Z3DW9NPExzm7PeynbnHE/
f2FV6mXxI/Z2JHWcSbewUudGOsvVUpO5yoWqGG0pfp5FT1A/wEtNQ+7/Z61EB6H5
ULBgvlyR7UMHCM6P8H5i9fZlGeYCFYMw3MQHYjX/didQQgNQvYiQfvN/NnsqFo1c
ZQAGAtUj0PQYKDIIAr7Gx84+cOBFcpdSDVe1Fv73wIiUYqA2dvJ1rnvd5jho+sYm
OM3ifxCyXu1DXn4kayMl2+WOu8T/5b8FRG3L/HjvG6TRtbYQFtGQs4jDoxuDBj/6
IlJeLZJkrptFCV81a0TGv2avZcN3L7n96/S06+ZmaUFdAO+s/WBbhkkdVQcsWGdi
IPlD8JHZho6FE/VckyejQdUbY5ROrrbRLdB+tntZEFh2TtBFs/qpI6R14AbZdJaw
VKV8LFkgzQJMaISoNQ0i7b2HbZfQQ+G7cTpzwswr9P/8AkWqvlO0R3UqfuhBp4Wk
Do4sMTDggiY52190x440FXJlq68Mr9MCWczdmSTZLUlLDM1WdU4hPUWEhEbhPLW8
wvhCBqsi2BzdRrCb38g/71gLZLcnJGO1fKS3mdiCYC53aLVCOGrCZ3zhDtcqMErg
TOhI+9eKu+2HYuAjHKnNKgAf5K2wLsu/Krw/waXtRBNzEJ8EV4zeKONsCQbfsdgR
B7i6CCspeBSAI25pDJGv99SDG0nOSGrGB3EspJjD8JL3ZVP6LE7KvBiVqcMuB8uS
orQzAYGGm2VCH7rvvSEv4rn8Tng6s60oC3okEtlLijFWyuSdLvCDiTNztq6R+ADC
DPKK/TeZCYRHRsiWqHP8gLx7cxCgjyOgNVqaauKbmHz2R6LPiWGPPFyeFY4cyc3E
TmK8BapBz0R6BWcg9bU8X2bLoRosf64F1Qza1KTUaL+EQ4HvuxMnbU1UawosPsV9
DRYwp6GtoT/r2NhBh8K8xztJqiqiN1iFP6V3+e07ZvorxLCQCRAdmUk3g+ZWzejT
cdcVFosgTG5OSe5ymriu8f/Fn2h8hDAdT3ePcjNkw8hahyDGcKXw2Z3J3BHqU7DE
edMZd4/b+Hy6I0q3pL6ssngHlX+jdZcP5ATbkOTFZMjJLkw4XG4R2E+VujdxISwl
vGpYPm4xZgYp+/7lkrCSdRWzf743SvXC2DbwdNIabDHCy4GdMndgDBvOs3VAImyg
/Vktn1RUeq+SG3uZ/PkFqCoW7rfV/Cj9KrRZ8IXiKSyJjZgRPhibhLUMnp7Ts3K/
J5EnWs2lG0CKadpFBgVgG43kbbuuPpo2L1K0zFMqx087fmpnBx2qdvBvXrA6M+c2
Z0NOEqYFpm0LIWUtU3Kcn9Adi3JgrBoZtJ10fu0JUWwzdDBPAHVVkkJ9CZHyE2mZ
GGCeMGknNFwUFZu/lmIUeVSlFtqSnHsvO6hWeFWcdtNTN/CPEieyzBg3mH3NVNJD
30ZI3SnwVry+ThW025YsdIK4XiqZuFt10KEjwves0WEAJeGaa9SGKU4Tcmcxm7yf
iAb3mh34961SrnOnwVxomfT9xx2t/aVFT0GIOr2GyZxZKac3w88syMwfn1PlhjvP
2gbaPzeoK41j+E8k13kkkymqGAsogNJxgxT2FwqWuGMuOBJ7yXl++jFBQpBDFIzf
bUnbR3ArwTZpcXANi+Sx4jX6rKaHd+Il6V6CTYNqLiXpgzWRqcHUVs5sgTjx+6/a
JqzMrjjLvR3D92rwTyfWyFH/bHARn4xvAEtayR2z2Btr2hfzj/VIFdlHwPo1zVEx
McFyHze6A+Owg2iVp8vjZKXYDVETcu9/m8B4KLjBXzcpr7HVxBbu0ZKUG1jROQ1N
8dCVRycMeCoLZ3sj8VI8Q77ZS+EvW7g+RQ2ZipyWjGKVP/D0hjnx5ggbbKAyX9my
Sv2w4dKEULwHwSC7MWQZcTSwPxMDeOkOE08p+lYpakJ8Rzep/DuYEXvRCfBciUap
N3TmZD9POAL82xQY2jmKMIS7KUxco1vb1mnDVvf8OJoyb3vMYXVnJH8GwvA9Qv8Z
KZyrHNgIP5zbmDHKBaKcpw9sU7XC4hyJZkF/dqfkgueMPQ8HhMYBoTIPSdQyEnJX
pS9yW2YwtGb4Udku7XhANdhJPETwFqxysq6NKmcFcb0B0I213VHnT4MNtAMojfUr
dDXGzYrqgkGAyiuWUKExQZ7Lftp31kRfxJFQh+D+py8vgFApY43GLP91K3TR1gPk
MiXvVvMK6ReMCiuxX+h/kRhFUTtcjBrI/8r8CeZxdr6m+YK5rO6pOr7CKtNaF89s
kgDIxox9qQARioIVr6/fcp0JgUiML1FzODWS45tawoa5AVVsnm51eQKnqImMSVLq
E60hrwEfy+SfHtp4Vp5xsMGhZQG6t0s2aNSYess0H65r54FfRk7iVNL1QORFIjFS
SaqMloKeBF1yFpwuTw7cVx7Jzmm8Y2I9M+VTi66tv0oIBijS9CpfVRx30p+TIOiD
L9yzeEMI31RDDskeMt4s6G/fWH/Xr9PbVBNWSOprR8LKzwZ40XXXSE0noujtO4Yn
uLXye3HK+9xbxxkCyorHKZSZVptsF5dCtHnOMkBptZbHsPAvIp7GsU4Sx4X2FDZw
R4MXDlNk0mHCxPbGBNAw6mly2H8OzTyltVez4ajdAesf27T1lyqojnBQCSj7oXKd
sgc8Svk+ARC1mfqj/PSaEKrfGqKFsttSCiDcdwjuMP3zKugh0Xveo1RZHpTIyTAT
r3sbSNty1KtqUNDkAB5O8pIq4EdMfofXpcUxPHtTjaFFfVGutqalV3sX0RwufW86
ShtMyvrQZRRwmukvFQX/+2XsJF88PrEpxWmPBhxWSYwg741O3tL9GocEnvV3MiNi
EwRYYHJXtdZTLJGMgibZcjY4RMgF/Hh+Xxg9Rnc2bB9j38xXgP1vFSEsvRmdOeba
BItrY9TK/BzwXhYve5AAHZ+lfnbryq0YOU+MKh5M3dLWYjHaxpw6y4+parKpib1Z
uqInZTlFdi+VzCx4/JC+ABBrSvHUJnMYYXW3idMpEqngA8wZxy6QwsMmqgy12Jfl
OuJh7jOY5jeArPlYOFigaPgVqy3IxOcurVR3YvWUBtUJvrmrxWxtEFKtMo6gMwV/
OX4sPM+syUu63aty6ioIkZwKWMXv/a7VI1vV/LgnxwNWkQllCNB8btrjQfZlkuQx
UiMh4EUvTbJ9NmxdsQ3eBuzWzi2ScVFo5R20RNd9hw41/gvnHv6Rl7yxAIf44b+b
Je/r1AY/mPnHcYf6taPSD5pJ6aIBPmXVSsHtZ79AXi9MWttWnL9wBJpizkK5zi+e
jZJYoDHL0YJRKYbaSvsZS0DRbclHnnFNgWWNK1Idqh2+2a5pT3OOoj/U7dvWk+5Q
QSrxmJRCaFhr/7KAGEf3WIXVcpP5Ga0FfUm6vMVN63SwVdfbeFKPAUUwNTogcf0m
TzywoJaz1ZRa3Ja1cJ+tPII4e4DFIMQnZw3mrUVpxaC0D1zM1lunXPeNJW9zLhHm
U0hn36QD/PyWd01yHYIwxTIJ6du588nktmjIGaAX/rIphyOVOtPSYcP06pvdUUL+
X2CB/k6CZGjLY0KGOJxJ9jQM57DNI3WzRm1Z2Oo/88FeakH5+KwfbqRlSA227GCX
IxCZgl46YZWEUTEw1FAItvKdjVpvxeyO4M9ih/OWgqvivlYGABjgfqVTiUGkWNBO
7eH1/pOlovrwKAIj4JLPDAsDSTlna5dbrWdiyKjaNpiyWbJG2yduGodIUpMoq+K2
4d/E9FXT0VpxN27JnVOcfdaLJ0qYZyojljB293uPhqEKERpuls35e9VjwbcfKHnj
Fd+pPCbPanESVvv044Ixm3/pwINgscuOf/tmSuKqzFnxQJCJM+Szw66ptPPccjEr
lpge3K+x+j8d+dnLB34zPmyg22aG1MHg10Lu9mOnKhZ9y3zsUYx8ylEZMWbSTIOc
M6gw1R1t8mduN1CRmgdU6sMTS0cmeYlRDn5+/5stYo3ZQ/XLldWDxtU7lJ9QtxjS
mAdRAuxr5q6o4gTdyjn24pkEImhw+aXQM0xuanCO8wNzDOsC+plRNLbGZILhAl6E
9yzjKMasPqFvZGvJ4jzhuWhTNEtHkWMrqe4svTxm4CgiEM5zgKg0RGc7fEaVkufd
c4KYdnRCV37ZZzTHpbBLMSNwOFb+kR0peUqOt0WhkXrvZAKxfyW5FG6eWPKv9xa+
12M7mQOdP5vM96/wlhNmGd0S/z0cFro0nBhxXxrFn0ouEBI14Pf+emSunwSzueQ5
8A4ICyFy07p5aoWlNkoTczDBedFC1Y1MIQdILePSCZPZEOvzG7D17JecYnV7dPtD
E6shX8y/mMEHndss+fnu4VtA8er4dV8TEKN4aZ9KbQJhHju7FSyZheNZVq6wOqK+
282rZtWysWfkqAYkL/QmwU2OvgCXz3WnDbvY9lmFzMpOCh/uDAvplmL+8iQPelDQ
gvzI/USHefLnAike958/zcw2kOVwTdY4iITZyAxcvA0E6zg9Tpye2x1fcJ3zMOAn
gW48unBveFc++9hxLLeDMe65AITR4CkCfmr9ooHhlp7pbJeh7+nT4IGBfK/EmSHH
M8bHUlNcYMzCahMP1XszdxEoHqCTahElgb4KxQOVAUTTXOiDMq26emU6VjZeX1At
xVZlv/SWydm+7Uj4N/KFyZLOUEvjsMi0h2RZ3EKzT7t2L0EQnWfeQaGxindW2wWu
LJGc3eo8ySDWbifeMxdiarEZ0KBCdkC0OwNwr22wle/ELcEDU1mhlfMrTHhkIvcs
IR7WwdZnE9iBi+j7+iWfdn4FKdZMOtQ11VIqMa3c4gx1IBOCRZpheOACqhTI95rz
bdZlf6OvxvsbgvKOIhR+23ShKRmJUuJl2SXhga1hR4XcdTc4+gRUfJdZRLIl6b3/
tY9W6nCG54wcyHvyjJU9Z4QfE2PvL6PdNjkVZTPmQf0XZMdWcw9ya9I4QZxDkfCv
+uXTBSrp2RKmlmAy9E9EO3vZyl63wgd76OGQrOa5K1PfaUScUlDhs7cM/mJDUq9z
J0NizlYhLJ+AdQeymjVByNoSBJxISAftInZtBqwMUW8tjK/aQqCloub2pGP+BtWx
dzRxwxrbz1NaFTivz+Ej1d7Zd/aDEP4UjrpfC8NEz69/C3YNNqFYkwkPUuEuMkcE
yqsHRtt9QtyHgVHJWqTwUqP1yYIX0P03gfcHL/vMk2mwsIC1gSLbakQYFThQy8Gu
aZNyjokXRZd0Bcv1F2gMfkMYZh5whG2Ryc5Y3mSe9Gms2ksiWFzygbezYJZZucXG
e693LTcvdQ8Pd3wmRNWaLxWL2JlUTqg2Km6mXLdRWVYU+Po7dRmY+m4tJz7bynjw
P3JEpkgiz7lVlP9qVpKAqblgywRREq4ud54Hk1sWziST1ZLMsIVc7gtCBWNjgLDx
eHqCbeqo+jcfnEUwrEWguCm7dFnAYIjwZDm2UV290UK/KhEUZ8e+l40/4u940fui
asGlsWW1Gw8lurxfwZYXUXqSJdD856hNfQuObhXMCQwM4smIWvyFoUfh9Y3vZU4b
F15TzIZdMqtIf2A7EgD50jSXeyz0xzJ1LAIWaHM26aB7lcTGnvRnx5VMaO3kihMt
xXVb65Uhl3DIQ2LI3VWECkuBAuu/zsTEvx/ZukzZ76EZGvKCQ8SXWAQoorE3VIX7
SL2Rt3vz5R0yOPFuiJlHEdt4S++/Sngt372wX1eg+CzWOf6+hDtmza4+L3m2cKng
xMOAo2oAixGR+kLYeb4+3oyMIdSURvv1klr0UCHqf3Js2oFyDOKMBB9TMhgFAIQH
rDxmvU/Bwt6zihCDAJFm/2ZCFUTj7iGgftCukTjNRRcwLC2C5owrhYyns0GAr9rU
tcsCaMcB2vBqJAJk9iu1obX+NsoLMMtvpb3aXugPsSJVqAobpAxrreFjkSCQfqTW
GqjoelvjBqOnuskQ5F1QImiGyxwOYTvvoaRJiWf2pNF7AkDVtMXJMEuWPNwvYXgM
PIQXDVWfxx5lS4MQpgkiHHYIVJVCUCmIyHqEvLh92qWKAhxCMv2raIjUSQ3ohW5Y
z+LlMECq9Tpr/iOnXp2jqAm5mzPwZvQBnhZrUIQZpK52Wxv9a7SesMNTfljf/ouH
wrfzUNfJW6Xzkiyl1/i1w/jjfhyOYq7ZStheQf5fSobKaEFv8N2UUDJKDZf6fwas
ne5rbXdjHB5qGmd8iNdQRqWfkgb/twW1NRc97s9gDvyX9D24wQ6TeacEzxh831JG
vLNwFgSUyZL6zwmPmDtY8FVFZB00ZHl85VVqufjDsQchkxQdQjVFzY+rc1Fqa5ju
sfafO93M6wI09xIF/gcPuKQdDJSnVm5cOAhG4XLNqSG58Neqmh7Dm8FXgbCJihuH
+ADY0F73ALRJ5HurIAviX2tjZ3txnx8HAY2/qPI6v+ZfXcbOTGizKdrkk3sGG7pY
+mbAqH+226do0F9Ctl/q1E2KpGJBPmIqFTtoxc8qAuYaBvrCq9ha+aCvAEgbo2jS
L/GE+jDXH+3XEJQCdgT2LGZJeuwpgBDdkRV8fOepFhW647DgWyKI2wu7HoLtgqht
hNUJQTYbLN2qcRUTaHkyDV+4EcwKqCqxpjqgbn1+0SxpC4kzKk1wlF3y5y/nCZ4O
P59rMPdd2nLjEgr5JuIlib/NW6zE4nq9/HtaInm4Copv0824HLZfkiwx7RGRmeag
0jIwNqLtaSwG5nUgOHJDcePdt+VcO+RxESz2+73M/2qZY6MUjr8yGsNZ1CkuulZV
T2ggkz9ZsAKLFnmRTUzkGsdM1PjvQsJxzHXTNj9hD+JgE6Pi41Ywuua55MG0O99T
QzD8vEZf9cRIxUCS74XL6zzYf3p4/i0N8TK6Eidrk80+xnXYORxJbIIBAWJimzqo
QsV7whnSUjPmO+jRb8op0BLxbZrXGDPnZFLFutlCiXQIHi0eG5KZjCc2J+Q/loZv
EEGmPIWS2YmeabDNVKInTmoTj1RpFFflWbGKyTvUoYmEa8gI286sFGorcdjMj/ts
y/4ZYY8o3oa77rC/iT7OKKTlQIyKrpfjdxzKUPWT3/9dSlurZHTnmAY5sCPxEv/W
equnqnLvZ6WLTarfblYDp/EySMlVeMAqCv9/z6Zkku1YJ1MaK4SO/YLqvXoZ1wyo
BTNoGmlUyCOgEYVhWjxymiB7QuvEsW+bXJ+tOsibje2RvkxTTOTwnEV5JYxFWLDR
lINdJs8G3WPmoeUKMu37Bqh8RSaE/d8yUHYjBYB0+mACBSK+IiMy549yGI5fLc8p
MOz+k2fDCFPhzwx64clsUpuwbymP2JGZ1vGbk9w1eeKi1Rx7WXtznm2/fTnxhnig
FKFeI5VSIWBKmAshdooRlfGHBfZBMtQSJcHC10QgH+lz/nhC9zhuUU7T8rpJyDXS
lxmeFaLOHwcW7EziGRG6c/uqs7JSDiq2SSDTdwco/YnAL8WNrOhyltut7ZP6DoAU
sqhjjwgPpl10BR8WozhnoajRPZDEJL80VFgSKOuQgyPDQrnMvcZXWyn7Ty7SXWXm
djy6980YRhbG93jpCy8RBCvvB812uXiltINW9dZpu+vDDRRN04qoF53GCTPyYTvX
rfKrRZPiHy+oTIcBuyvxy3z4rwxeuTijsxABt7UDRGRYU7bY3w6cimFFOopDUYsX
x8bYX6HzMMds1K0FMwxYI6atIGpzwAk+ahnoo/R0sH3Zpn+JJvHn5c0MtWtvV6Lo
cjHv37eltBWtRJXfq8doyUEEBQqbqK60FxVsqXpZ0J17/qXz3yb/qoajT6CmVOvq
iQ44UXT9wkMDL2D5eRHJvqy7X/KJ6xZyH6ud6JuQVZqKLop6Mz0Qg+upWufdvk92
gZtLo5/kyIjutgtStNlDRJ8M5s/LZJeIHSpXA5i+VrPdnQla4maR5r6C1cb36XE4
sqiNZ9F+CqqZuByz2Rk8nk2B6Apmw12kqhWLxGU9leSbYTauQexsbJpgiVdjcGXJ
UcMtj6rXL4keiPnA+6DnGKnSEg/pyd/MowaZW2KBCtAkntqC2KHtQ1+H6Py4W4mL
vlmIQ3t3C2hfbA6nsx0/ZztX9WEEb7/61bZe2VUFPqc0CgyJUr3kzA9oAvfcl65a
rz89iLBNuvrVaWFMC3u/7Yq3E5JrRSVTB4tIku2OHuBIITXK02hkEtSH40icKTex
k1S58Bp6dPi/DEq6dKVDG/2p6TsAUogJDDEUztdi5pwGdxs5qd+6KMdLdGVG4Ev/
SF/0XgGRIRA7hfkUkVUIDRJPuTJHS+p95tT6tr+freL+GJ2WZOW8q3gDy7NtpNN8
SKwBjMwOTSTCP6Lz1JWdGjWueAVm0W9vH4LwgHaSs6qZfCU9sq1zAOufxPcRwzTR
AZHnHOVLtv/KEbhPUm3LJ5k6CLovfiBkf0AgW0WW66l3b+fgAeAv6nu+PiaIGZRa
bfS128UiRPFDmqk+8d9LLJ47kuDEYacyRZpVAkboFtZR29bCe4qlQ5g9XB0ZdouN
gGZJFNmLYZap0oXyTEsJkbNEjqMa0RzAU+BIIbsdNsUFYayPal1/tFvVKqvHKMdi
Wpne3bdaxHdRF+MTqe9luRwRhDPMmV1tVbjlPnb41G0/8uGYBvJTJ2jJhWLcdSjl
atePpnNWXiUa2UO7E2AH7gxjjtIby1rK0jlIftmcOTg9dqOHVMRt0Rg52nSJ+slI
58IK04bKVKSEfWlMd5tmbsVdBdnNXPy4ByBTuaoXw9vEUc1m3BCSGubkmrqjCVpN
P/aoUDKDeeJtzSZ38seGb9hCPgVoAwyMz1mF6cTvH3rMezKmA4BXe/mtbJguiSJA
B4iosMan+ZjPOX1X6u0QSf2oa4XhCiMttxCZz1vNCtbSNu02H0pfZU0u4jA0uD41
3U3uSadLCc/oP4aUELzZnRw4pB6wZLJi2vr55806XO5MxuKxaaLApsev3YB2c9G1
xIBjKE6slkbz2bG5nTKDv5j0UCqvL2jZ0214j4CJB8euMuukTK/kVGS2GkQwHX9k
YUvPwRi3mFkGYWHShnRiOEszabFwnUdGkEDW8tWkONyp/qjke57KHxcCHwA8fjRh
57y5dxcNeqA3gGOuTyRKynAmcd2GAOAXhEFfzW9s7THqU+qD2uPmof7YSTO4Dx1j
DPgx56l5zqlDlslIq4WrIUvAN4qXnknrQA/IjpmFx1pmo7ueV1r8aJ3GaymGh5zI
eu3GNKoHWuQYaG35++mIH8gdBGpQN2i440hRe8jyeAzDN8e/55w8KFi4oxFcbBl0
mtxWEwm7rG/19jo76OZth6N14ojuZ7lP9+OWOKuzFoYObk5whxOGD1YqMUia7w0y
Tw30i/ewnNi7R5wBr9i6CAyV+DWzfM5dcMpI3XaxXvbwggcmbrv1c4h2OqhQAgVi
Fo0NBTKv7m2khfd4mqRN3RvRjv9/u5/B8tBpmvYg1Wd9C6O8cAdfoTVIXFxhhERO
lLLEOwdXiv9V0C+meKWIrQJAcXFOZg3fl3/I7R0qQ1GELrdx+wcxbFId5JTo7qAp
g3ftVTlj7U7P44JVaH5EWDdIZwCLwFyMaBXd9pzdLvw9qeI7hAg2MXcyFqy398gU
Z2OoTw1IByTzDDckecw1b+lLG98PhK8nm0+AIsEtKHC6F39SNK2CpOFM91vGWG7f
Ultvs+LurMYwEMIvyCrBtHsVZo2Y7YywmGzG4p0pcj8QjmGsDxbuL4C6upfwJgZI
RLzZ3+XDm2kRkVYG5U16sMhXpNN0/pED4ooA6ob0Vt8G0/fAVQ9FLTLj0nNFPr/k
Wu1xewV3Tu9SyM5Xedc8yn3yHIkcJivpfiX4LOhuMRiTlG4DSzcbkSdPMyRrnc7z
pZo1RO2BLtm3Lhtxmh3vS0vkn77Bj+beeSgoRk0vd1vAEpQn2nFt4i/HNT/twLDM
LkBMbplXvak0hYHPE3SViGLTNRfxMv88girQrDuWy5XQHrL3LlnIfkra/5rShrK0
ClaTYIyk1AtYWch0HHMn6iUKQZgdn/R93q4T44qRSaOZseNV+bZ5vgTaDT27cZ59
wdCjxRZ5N6rIM07KHUPYNqmhplEa2dFzFbtta/wH/7EApZmW1WZS5vY42qpnJBxv
ks6IU+Gb/ZgOdUhRkhv6K4zxYIwrTOJ22Qg2obPb+d3okaZkHT+zrR75g5PMWz6z
EiPg2ATTEDDGvIVpv/AwKXuqDDjzz4qAJB5ryfb6lA67/IbO8qSdkmU2dVNM8/0o
nOnI6heUjnfeYq2jsxq/N4fwx/+P9IV3QYasoF+qe+KMiaY4W0oJwh5WHeV57SMP
tXEIXaGBcZzEibFFK9Dw2cZyo+SveqGocMu0WDKDl/CRki6KJmwKTvCaMRhbnL/O
+RzBzLGdFgg39zXlTtYtJsjrwjI8RDmNX1y7QFDFAKsn6Md8Uwn6svd2mIMXk/Ww
Y3xvOMJBt7a/6JAmQL6gnWi76rO9CsyoCxkJxVL+oSvQtjAXHxyvfFDBf1K5GDaR
4cuH5I0n75HCWP0czm4aT0ZvMU44iLoDGo+OcXTHZ22sy6G6uW0lsQhG9p5/JwcE
8TxCKFzDlA2XC2BBw6ZApOgzDg9RtINbUwPitNYVigrBI+S1zPUc3UUJEONTDqlm
cxRpdsRK/nzudAehNe8yYSnYOVdRpmAcVW7y+gcF9XdmDbV0DxE02xuqIfQupLfc
pRtrmlLI8+NmyUr/D5g+Cp6CS/S1xdHIO4gDOtYtA9LVyeF6xuMjbbX+Jn2sUgUh
XjyFY53DmNqULC2cAuTDtLDge9iiwtVRFSdW7DKk0VpO9SaCl+8QnqEJfqBKSUnn
n9dRQR5yThE9m5a//eT4AG7xUXpRIaykLXnnS9ckyrzsAqy4+XNV9NgKniXXTpBr
MY84dDCGnuuoR+IsqU+VQF2w+VxQvztqZiKeLi07tKSv060rYs0t28jXjDHQw0W4
WF3pOop55rg63G3B/NaHuOdFL6tCc4ldhTlUd9TJ4XrsZ3h8TIFw3Nj4p9Blncej
J7t4r5TdHzjayJX8TyetI9xQpWToqro0BqDaly2s1lb9/jI4pdKHb23afMkFIN+e
VhAFuoQemeNKU6YDa3BJ5nwehDXw0QVTWpc9Whk1ZxNw6EsL7WSkFv7a+ou6cVya
sVtZbA70UVbwHjMF1QxWD2Twhpd0AGwB5FruRyH4Yp1xVut7fK+r2oRWsRAJW9zA
zEpdP8Lwa9sWEsXjU3DIJNQV4XT1VzHNVQbJ0vUHu7Y=
`pragma protect end_protected
