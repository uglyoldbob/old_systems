--
--Written by GowinSynthesis
--Tool Version "V1.9.9.03 Education"
--Tue Nov 26 15:29:30 2024

--Source file index table:
--file0 "\/home/thomas/old_systems/nes/hdl/temp/FIFO/fifo_define.v"
--file1 "\/home/thomas/old_systems/nes/hdl/temp/FIFO/fifo_parameter.v"
--file2 "\/home/thomas/gowin/IDE/ipcore/FIFO/data/edc.v"
--file3 "\/home/thomas/gowin/IDE/ipcore/FIFO/data/fifo.v"
--file4 "\/home/thomas/gowin/IDE/ipcore/FIFO/data/fifo_top.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
bM/DxQX8bp/+HIoZVMOChzkokrxQxW95yKsZpJKGxCMidk5mOAraeH8JZ3AAZO4E5UX9mzIm4i7L
a6OJVNT8KZDy6UYf1HNz+nsP9CztOAAxf0XiY3C4Na2DXCaE2GuQsNVpgk9wekJVrqblSAXKOuOT
+Zbv+sYqx7DkUJhqSbOG16j4xoz9V7HotwaLcP9x9D0xITlflARwxmXsej+N+Ud+K0epu6BgFVSE
nG8OXS+KmIPpK3yCpn7avYou3xFK7Jg5dGWaLfNuTlORx8e+qNSJLRfvq6/SCFdzHf5V0kOkNcUS
YP8ZLam+mK+7zxuPY+/OA+2nwURjZKkZIYW5Xg==

`protect encoding=(enctype="base64", line_length=76, bytes=139344)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
fpP3RLeqg3wyqoX8c+mV3s28lBQBovH0ft6/3GOp0zHzkyVPn/sZQSqk0UH7UmsdOLc/dGfVlBwk
MKEvoqhtvFdJZpk+fqsGCTSXnTcka6yHsUTrJtaoTRc/2z1b76ELde+TJRwJ7TKIDKhQK7cymsWv
kmMmbQGBGtUWz20HWEY39T1fgwmI0YAX592sOeHcJJSiI7hfZd6+Llh6fXtPqwlz8RWbTMP3XyhZ
BMjx9Cyc1aePhGnmoYohLg0tzwQiTN3wJL47jbS6wStgiwkvM1tqq+KkgEsLzA2NEj8MmKzLYwFt
q2GtsOgwVKTtm2VMF3Ercrz733SbJTY+LNKhMakmnBVjfb9GryFXpPPAX+rNE505SbV50nZKOvVN
IXm/zSVWDsa3arXuoDZILqYqrwPKMybYRvLul/3isn7VXDRa5ghwP3tsNY5QgQPy8hk6ttFCXHcy
fukBY2Wy5cR4kBS1vfwWEad8rhqNQIi+j7W+ewz93QYjO6nxdZNdu+cuYJKcXDrDqXj7SUno+pqq
CzMfu0NnzWr2Q5VaYUopjsVJiUtPom6PcKKpYH8mKbrDffAu38GGOwAKc+5GVZ/0Dp+SEYdxUvWe
BoIdmJEdyYOqLq7Qna0T853JARRL7ZiusgbmG4SSAieDUB3cNRvfuPAnyDSNnBVkc/F3gGSNoEmp
/ok8cm7X/ViMwEn36S9IOFdFqFQSI/4vA0rMr4b42l61Htc7cCkx04VvBjPNh07sF2Q6sn604dsK
upefVcgfNqN48Myv6OXgAB9Spp1RkoFk1fgoRVgEO746jNZdymqh09chrjZq2zw0sd9idvVTgkxB
BvSoV+uLgZZoUQQOimDJbA8uTkmOD7SLCJt3QTjhXDZTcH5th2p2N7QnZFlRKl5ZwBhlCKytzlMv
Q+gVp7EBn0Id+ne3lyVN6cn2lWR/n9UZ80raBUB4Y8qpZK1wc5RRSiQlcRuirLXKCiViwOmsrzse
BC9JGrT/5SFth1X9UwQumlxDZvapy5LBvTMtk5nXUqxO4IovcJb28I9kGaCb71ePAf/2+mAdX0iy
/os48IrVcL3UsrfXP2FQzMHkVpWBOXXtC4NEMCAOL7+0ZDfg9k9lFlfm7I5co5mFwOOyJL8sdq7v
6V2IaDZ9QKzZDvYxjjC3ld19H0dPapEB0kpILwB/WqTnRyIAYCeeIbyPILhkkHiQTOptE8d/cOq5
hJTdTO0buBWsFk6ktudBLZqbFSirlNcZ8eD5296VCmzzJD0HxnoU/tKJ5i5ES8pruuEcAWVYdrQb
70KhSwd5vuzOFSTbY38ZyrKg/1+t+Dz+HX35rbs7/B90g6Y6oC6WFc+mQlU0HVF+7A4HY7C9mkLT
bS2IPqSeVwVSYYWipQt5zD+oUtMFfbP03+4aTeepZ3XAAU/eQ8Jx0lNJ4Bu7kW/HVvyS8uDMqLKs
Y5N4qLu3VTXhR0O5wsKKNrQQkeo0SoeOAoTYe2pWk9wdFGsT519w9kTKh7MaVn+uu013FfiZEybG
FQizKx5ngyA5LAbhFTQoRu8gku0Yqwo0Pkb5CGWs+4njkMpPwLgZbV+Hf9Yx0iKz8qrA22teriK0
Vsajv1kmVLSnuuz3UqleKXJnS0KaEu6leGecmpDuqCXpq5Y1N4XoZTuCkOkcKSLvwhQuBhieIX/0
uRYAzjWt0V3CjvKx4Nn2o07GyMl8BKdeK842ZCNKD/SpetDLPs0WIJiOZA8WXiq42s7i/1TE0CL+
yON9nOwfNF7KNlCmucveHjWM9Lb93UPR2fBspnoRbfi+b3Pk+qHCK6/kdC3RC4EGrduUHuHEIpFt
kpLxjDNrT+n4WajVpJ+u8G4ndd6x/9bL2Wu2GZBvZQ+G2nxZjQXM45ZkAbDyZtcAm0nVHa9rnYle
vh8GgD0LbzWW3mVAJxUoUSdmjnWzplkmol7rzHJgkrq2LNUvewVZJR+bx+Gi0QJvHn5WsXMBKPjm
DTSK+lwLqoyfTS3HdLl4z/Bitv82Rf870s7eVbtSWyQE5cyurRya3uEFuiUQjXm+HArN78qzsNfE
lbJ4agDikPI7twQk/25YVPNMDQNUydaA4w3xBObJjihyv0iLDt0fICe92gQedRQ4nu+4zrNIVgv8
qQX43n13TmyQ/jsheQpgykuvP1n1JZmJM2hdNciCO4qVCey+/DkjfClCjwjj81aE/Lkmu3/mIxUB
YAECznMDHVj+O9/Z6Ony2s9Jm/gn9jxzQGhUxNzepr9E5jHRKnGm0CCgEKjPzGz+OcwgJjuluLYd
0HXUldRuSukUkUkGs/YNbKF7MfOpoubzrggdoA2g/kom+yoyGSWKPCD8GYs2vGjHvFwHTiSwu6QF
XzVIFpat1LeC/Rwm17G3+Sh7hBehAXU1LQmkStzfxG2MYnuMLjhdpzZ8vYh8o/urxXcE6TpVTMA8
ugMX6InkPgPBKZlCewdb/NelXzphmp862Gacek35ouhNwZfqJMWAYwnKV7hP6aEPICak+C4rJE8I
1tS1puS1BXSvT0xfJ8ApwhXGdtNSgLVmxu7+1rjeRXkp6z7hIDitkmfeMNONiHHuvN6RvQpoyZIW
8sE8UhVdpWmL97hUkac3k8eId6WypmVVUoiegiVBNzKWh5+raqMRoNs3mwAwS5/HIpZRRIGfkPvY
bKHSmWAfc70kCVN7bBwQ/rwM8e8axZcKP9JgQKaSCs30JDUqI+n6CknxR3DI1psNqkgf2ftkQkFK
lDL+LN8OAnldnlYMQb2RcYLD9y/YgdH+Mb4th4DZxleFjqO8paFk5wxKg45fVTdkzu3nZbsg2Bqq
K2lYRWXQHKBtlVYJ0Ag/Xms+RfFZQnKJVwGyPgWYg4ZDH8fgypU0a9TvhGYopSLeymWPLWDVrSj4
yrEZhXiC/56NiC5Iy0DbzFC5zcOlhKjDXZdYwGZ4wlv7M0HaEEWv4ChSXUGbvtuemGK4D/OEFYCm
VlvYDzNQCRHfkXK8zRnstaqVwD9d9WbWg8qTnLNPuCLe20L0PLubYfDaISeh8bz7/QAjm2QZxG5n
wbSd0WYFkC2++5F9xuV7IlTXEOA72NCc4l+egGaaYHLYOMArGIyEFsiwrtlCGf+t1dECOkufXiIo
m0gPxjDLiDFptWiDZHJhf80HMSswjWp3A5iBRGg1vqz1tzgmfrnFgWWqjS6U2tXwJouTbgvkru3L
5FJPKVb0edf9lXl8eIjccKHt5kdFvo1AqvSLswZf1f1R6AeEm5g0KFdqueeBoZX5quTrgYL+nNGC
n1gdXztdK44DeLt7BaBUsF7nOk3qZs8JTuZ2DfL9Ub8jer/xArfxFkpGNpRrQnKWfF9vlG6BCZ7G
BDu37dFRwy+Fg0e+WM5VVxLP/IKnSlR5GTnWKXuZxX7z28I9VJiunVMQU8SchntfGPgPgAGK1d70
w1we0shUwBpSRh5NFjfarLQ+Kp61GfnwBcjDNn8LLLaMwa6n3mFniUZFgywHIKk4j5uy5Ll//FD3
wlH8g2KmgGtcH9Axx4TF+YA3sT+LdCaQBpRGvQm8vHMNn3XjObKTUGwUmR8YI6WSpZC5ok4CFsTw
fzzhGH8+hNSr/QDyHA38q9dFvlPTNjKJFsgJ+NVEDPZDjNFrc8NXJ55jJBNEq0g4Q1FKMOVPjK8F
gx3h2OCTiy9ld5dG3AxspqxFd4dRhHKmlD0Rt0TckJZb+aifXE5zcVHBvR07wseLpvf7+/Q52Ggj
fkPART+Aiw99hnjGyMCGFaE6aEPV2Fy3Ld2E47gk7sLyB+DkL+RV3645pYQyjSn9lao8JLnTn9Bx
IL7td9UDC3mATHHm1/sO23cnItv2ftop+sVPNst0mxdJHk04bu5Bl1TK8RMBr3kZ/lXRbCaWGriZ
0K0ipXQa6tsfG7cwL3AB//XKE0Zl0Wg2pD99icb23YuYGJBp/GPF30om3nGmPALgdB5BpOfl+zwr
hhqZyhg8CjhQZ0OgrCgDaWP8BQjXjdeO0Id0qcNfHj5HmXBxTRH3VjDiEBKncvI9nwdqtEOFvMAs
JazLBMW2xGZ8Kc+uhdBD/6ZI9Y1UfvYBwcWEQn0K2VxrR3qhpB660QGFqnCLJuqOgBwhACvjI9Zl
bSAntqXulXFvjueAjOHPNU9h66cUdlXD1MsSyflXDEHfdXWV/rglUe3++ujfvW8qlIMOBsOk42o4
diJORY1gr1IPiCD2+dyn/TF/0ee4XnjzItajAa6HdMEV/uqqoKBVRAhlND8wQgKs2WqOKoJCetKw
fasSXZ7tYNcdKKdFdPBg6D5RpYqG12N7I1Fq61CNnJ75Y1xSRp9H4Ix9pGmgfdJt6gFX8nXygEN8
nhZd/vBZ70KUWKCLK1OXE9aPp2JnSQP5w3hoVFX/8z6a6GzZXwGe+7EE0juYoB3tfBY7l7cPAB1h
SRG7PUQx35DfzQ3DDOGGnF98dVnCkQSXuh+FTMDv+U/AcSi2wbdMu0yuTZFfGadmxilhZATAGn/M
zLwBXCwu5Qcz+og/BDTwKlA/p+VvB1JoiPlJnLLlpE6nuNjlZZxzAGIoN2VyNe0SupPFNmqeRcrO
BgPfk/DG1wLQVcZixjVS4k9DcpzdmeTIYcmlb27iI3X6IIWqKU9OGHAdhOoCiQTDiH/GXaJIQ5TN
/n0O+hA9XZTdHevcl4Wq9WF9+P1TJK1ghHbgjCTOZqV0BYZfyv4aSyXGgRMpPM6XOvLd/BG1q4cv
qyz46zeHeg0Kb/PftbwiXAMVGgb3qVqh/jiU9cjZ7zZgrxvpv220vIOdYafwpGAA0wmLbL3vtUz4
LfP6o+tT8Y0yfX1thoO8c/2FNotCD6dAXKkw55tqmenp/ucs5GsKHbLppCe+SwTg2+NqqJdXufAF
ryB+g/CEKd79GbgLcUkl8HjQkrtDT7D4NYnLdghc3Z5LGuRPfCLqorTJs1B2LfnAPYqXOIUpc+H9
RQCCI9WiaxEZJNb5KqVge8XtPyOyuAOc7X73/wCVyV1VgkBGsjB5lCZPuNYRBG3OAr0ciG+rlZMM
gBEoW4Us4d6xrlO1ubDjCn0ZGEMJ+4Mzb8/8Gl6xYdxPwNF/m/FNj3kihm3vLxDaEA2q6jQ1UgH9
C+PI27xDQWzv8YIT6wFOd37q6DTicCGnREXS46xSR1qWx9vCC8kOg3QQSa+riGyWckPSyDx3MHep
4lZ4tr8sw4VyYMbzRTxBWDwcc6JHNJcuTiF6QVaO5NKsuIt58p+JBm0+VnnoKtIa1e+0GLqH5ofB
BMKQKUFbwYd8Yd2g/RrOQRtuZtO0/izZGS+O70orsEIfYO8bOshEAIuXsTtnf7hCJznzxZqeqWrS
L4WT486+LKn/VoseNi+4Aom3dQLHJuZD9yP7DKXNunDM4v2meUS7Vbm0dzfXTsRl0Sp0Gaq95Tz/
AYav2X3MKSEUWBAh8jgdF7o3WFNk/xg36boR9fy7sCh268yzZ2qeX2djaIZWFwaBaJ1DMgBHiMLV
HQXx9z9KsJlBIG6kK/VzHsD8QvJAQHC70yxUJMLK3lspAkz3/4TD/dJU233i9/rJkovl2eIg2QKj
FXpB5B3n42y/fU7wlQtmu5QxR4BVybJZnUlcQHXIyPpPilkAW5y9ItVnzgBEvAKiv9cLxj1xVqe3
P4nYEz5gHEhuK/gY8X9RI7Iz8eNv7K3XRV4ZPVxlmsJakhOFLuE5JV5LD0xCrl+hZ9pO0Wvovap4
+SNzl3VbRhXDGx+a24wq8gt21SxWu+jkzJiU2tRAxHCIT3l1pVYcUlZgoCT+CuhxtpS40h+dd0iy
pS7uVVPQnicB1vQ494/X20pYZY+af3oN6PyGBati6fUhRX3GrRBB7+qIpfAgHoeumkALZDdl7p1x
MgDfuO0CqVnae4+/CDrgBhn8y7k0UgDD8DF79+Sjks+8D95JoUej4yafEF1WK+MSrpRzW0aAcqwz
P14N4o3p0rZjYp8RT+8z6BV9UuBoOFbDM9bqMmL3VZAaaMajtAn3TthgYVq//eg+GJ4g6tES2etb
VUonvv8d4jpuBUk7DJqi6rqAM0OaeHoBWUDM2Ltd7EfVAeGksboNrQoZmGJK5Q8gnhpsNcrHQZc5
5yHXOJCQgFUfiEhUWmDLphLCxsjs05slJofCHW/IZc6DVdWAEhlOeCt6e1LplcKTjG1XyaFuoBlf
q0DbBwvAX5MvnCDJo9iKe1NqQn2tPcw87MGEoM8wdF1JxulRG56u/K3d2LmEoVdLgDNq5oZqVD79
evotySlMUNkYRFMJpjwfN7bM5f/mcL6FbVU3klDDqWOZtCnth/PpYA4pAKa4cR499cPjfLSCMcUU
UYHX6Q4fePy25SrUojijy3ntvqcwPL7EOG5KJFNniv1l6z3jfUh2DmLorx+NLJ9H6oqSK3ckXAEM
yfi6M2oRhFTCYvqKM+QupMmnf7aMPYZq5oZWJs3ZLC+Ha7uQGo2mc79DHfGHGGFkxDfLuRgcSorl
p0fqe0UJNjKwfxAhm2KWGH3k/aD9nVUpLIQVFWj8PcLJZIQ3eCo508NKNZgoFvt2LX56s1nVz/AE
c0wvAdc8HomULtT3Cs16Q90/Oqkid9f662RWwl/hHc7MtMJm8jKQHJcJlCTtg8XaPWMwnqHbJ7BT
WWrv54ToSrO3MVY4uY2Gf0hob6lEb+5fgSTmxM5y8ZEgQJW3Fqc5eKMh8FCMHYzlRsT50A4JcLSC
BvPQJczwSVBENQ/u+6QnLnNtovdjYXl0bXDCBIXEkDlX+Pnt+6vy6FYM8j1pAfP+XLVUlHoAmgHU
fReIRswkoIdctt0xOpkgZmh3rNZS7ZpHyL6tqb3UNOx8ZaW2GfUreEmDd4Lzh5YX3Q3BrBWhATns
umbXXaBjmB/7+RCaD5EYMCzqkyMtRFh0X3h2HPLJTQ1dzFaT1q39AHzd15aqcoljKeH1i8ACRXaY
Kdun55lV2/tk5Kr7f2JSvV7cY4ZyFclFAXlCJFKzhpxoYWFVlut3d+SU1jgQp9jqIqxsykqsn7FY
f8tfznw2yceHhARywyGy3tTwiusQXO9oh4GksZ1J9SxkTADd6u6iFNrc+h5nyf6OAn2hxdQwQBQA
qeBn4uHeqs2B0UbBOK29+zhHkQuvSOZPlnNHpUrXPytGAkNJYx6lSdvHN4tKAADHiYrXSUdwnMLa
XamRyOnoy3E6oXl2GwFzDjc08Iswnbobfo5h+6UvZycx8wrpDyVI0yJusUh2ZLMoBBSu1lUiwF+R
XzN8WfaX37c6ax0+vNrV9ecIrxajCPIA4pqveWweobeWucfRGbVidw8qHLZBl9PCV1yFKQAqEY+k
nntE89Hsq0P+dTw94sSQ7GvrVnEy2o7PCBHCu17AbYJsT61aCi1BIT75i44sDGKpOUShL8FBu8jw
Moh6OkGH+K3MS/vzZVmzco1POWo6bf3ndtK+mYEe9653wua94WYUVotcVFcyG0AAJWy3m7LijMin
kpvROvX5bI+IgSAxKOWbJbZLKEegWBGPP0uzNy2xAx1clHXbCOAV85eEe6er7yROMmcOsMH5fPeh
zgVGIWiRr45Zw5rA2+y7VxSiB9cB/UM/fmrZlmCEyDWTasXB3VL0ladwwEdGz+qGw6sWwDsr8C7s
y/WNhrj1Hht1vM4dhEMk91biN3BqScGF9GlHEQwsY6yNdNdbOkJ+xUex4E6JrPM+/sYFcoGRb5bY
hCvReQUPSHdpEbf9xeTfxDEGIvc2BDBi8hRbCNfxsMNSWAylwlyfh5WablR66U+SjbRXD3FjeC8I
YxnAEArqdDjPy4o5PU0qBeHRBM3lcQikyiFlnciI47BBH6iBAd4pWsBey85HzBqzNRkm7UlabvXl
Rpqg2BcNqj0XkKqzaXwwMhEld8F/2YeexxhroHjTs9HizmFzVP/KtqVuVUY/dNA2RaWt4TMj4l/o
G8H0jRS8nqJ60UUcMgJ4kttGmu0tb1CZ2MS2S30loMf7MxQyKRiXyXVOR6pCVvbw9FaM3R3ohcr+
kHN5HanKVAOMD8wEN+sj4uh7oyns7BegXudLVgyhGOfsTnIzMnvdRrHBw2sbYku54n0XyJzkMoZZ
X4PvtHg53//du7wAGnfQOX36osm7Lj5HeOBISISnqS17v/YHgHTac+QDzGoEjhGnqOK0Ru5EqZ4i
btUyMgPpKXxJyZ2yuySg1ZrwSmNGRGHle4yyKqAeiYzK3utKr1mgxtpev+oHd6h7ArWVGUgQvrn6
hi6Hzc12zJjt4SoiGBMcoHF4UPRSuSb2A4Hi+YEW0y8jLKUQBO+ZkD+vS3Mnxk0W9wd9N5SXx3Qs
/nqxTIasNJFcMG2h7wwhNtAccD2hKuZG5JhBINgTErwEYf7iY//Gl2TlhGPOuZLkGT0p/tCal4rA
6zncnCe4hbP1lQOeOBvy3rPeywFcsXag6pb6KAGJ7ZzC1rD9Lj6+3ofWtzI8tqrEHV1+UE8tVglP
wabXae5qnF3mXnu/2C34XeL0HdVbcLkAr04T3B8147bmsml9C7NvwYhDrERn0+5dVmOLd5/h+gbF
xB/n/iEox6yOYv3Pe9SwiroYdf/+LhfKGnvckwgMrpACIxcIjwVJQgVr51iI2QdbpRlGSxJqm8Iu
AxaY97wlaTtQBDWfAB0ZyqIWpVeDOda8lF8VRjKodet3RLyF6hDoCLA1OHGt8dBN8+8WB+T5AagH
vfLE8r5WuHizPgN6+edW1lMlPMVs2U0Bhq7w3XHZnGMZ5aDmdvTBdzNNI4ltHLvB9NCi0/LGPOwI
3dCfCS7vZlpV8Y55nIwQCz6OT8Sk6/+/6ZVvM8Trs71YPlcomIbn6frUlWCLpZgR0aK7gKWPfw8t
uKh9lH95CwFCl6dZOS+vredLzds5V/YGGoyyrmxukD23s+K9TTsSyUdUJ0KquLtwKDKcHzZ4ygW5
a1sUfSEe8WOq26iK9/aWaclUUzBtHAJFY20sclHXbEUAoxLGQStTGWbGDtXOzRp+7gYIcs/ploCT
Fltz/d61vWC9Q5Ol92ci4yCi9AdlaRJ1m8OB5qsdjvw5hmos+g9ANIT3xNMPTu/Ti0O86+WTtzxG
oMs+3byoSnTSng7PyB6AsRcIhgnNAlMNCLw9Gsce9OQCi9hBx3YTrtzCRpPzP/BjUBwjd6EyB3gd
YcGMMOM2AsV+OwAQ9nEdCy6h0sGvixsgvzH88piyK1RAYxzuGqdenCAN+kjWZh210qTddmqrcnjh
wlNZewZgNYvtAyIsgdoQizjkSAogfYV6ZOaHHvoGomLon3r/z61jf2pjeVE1Biy4dF/XnILrfFLr
AHZT+0gRwzQKdfKfaNKpxPFX0X3cpFm8TBZolSBTOISr43+q6zvdtaCP+2G82tjNLCynDu5YMMwl
e2seo/V/WlzUKOTz94KhWda99nS3oVmBVx5wBW1yQTU6XumOQc03JNcyrB9uQh/YtCvlWAQ8hXQK
WoKgEThHKW7us8wfbYWWFdjai+IV7HJSyT7LjpqdJZKzHpJLWj6pioGXm2pYGeU5MEA7MZ8otx9/
shPt9zSpRyZlRVX6PHhk+ygJtMRQwNHjc0yRh3OG2V+hX6pi+7qndISssQBG1UTGHYiZtIOb8Enn
yw07xitKj88b+3IqvJYoTwAV9eY41lHv9ssv+evdiGNbplGH3kNHrTAZqEP9OPtbdWZZDsgwnT/G
G1+gwV0OUKe+T+YTQU9kKtaqX/ziVjGukKmzQtZONumdkh4wPM5gYyxzgZu3onyNYICeY76ZXEAi
UE8/8J8yRozcorlXXL1DGI5kNhE+3g3Qul1/+d8EVoeblH0McxLs3VoNh6ti3hUYUHxeozXMEBI0
fOdhTYq82PCBs745hdnStY92d342rRMQ6LnN+S/ItuaK3YFxa6lntyFS6cjAwZiH9dwsxhqGkdVA
prM7mMvln1obPGSOASC75vhXFhbHAqyQR8pEgTcJuis7qVSqZ+pQDx17qyhEuoNb54HbH1+Hfe9w
AW546p6tbyj6NRM41ucvGWEJO4AwZdA1a7KELwsharnVqejBxBRmo4lihNAamBZ7N6bejifCHm8Y
i/KQatDiTPJ73pBf7ALAICk/L/l3RMFlg6WwbGIDyUzsg6SBip/cHE1nWE2xbSv/zfhcvZDPdcku
Y1QKp8QHWaDAwf77eArYDnkaGHBeOJYwGYHe0NJ3dYwN4H+7/yuMGIIrJRxfFUbFX623NTkH3MUO
bhyqVKZcUNaaWbJoCvvqhmqjlow7qT/nXdf8A/UoHs+T24cWtBcU3MiO79Vh37x4V1IU0MKAkFN4
QUTaqojOvbG6MSeCmhYLbO95v61r9n6Zp4eLx52CeFmqhlJfLOTJ6bh/J5d6nU5n10rTmVM5Nh3Q
EJJVL1/Mhqhw5DySGgKsGt88yFC8V/GQbm7LTaohSacCFQ626KLTifi4Qf8svrrKXAX+ZVoST4tV
V8wIbaw2EzcACogoXNr3w6EBcGPYUUYW/5H+woPMgAgJJdnH4IqVqTePOF6zmxCvjb2+J7UsnmER
HoQINsPOIYl6MP/wEFarKD6QJq2ZiBZEJYRzyBv0J3EpIkF6GNr2l/E5CE4ivzmTu6LrQmvkDkiB
y2mx2GdwcqCLxEwTFIK21HVeaKQpymxtLTnLtFczuyELPg1PD3v4iU2N812xbM1QHtlh3yAUZym7
ZWz0rsNV4/zD3+4hosgjfhWfiKOX1zFP0T8tv+i8MnRrbMnSgTSeMyEsqUjdkIp4kJOyQXT+Xgb5
gjXa4ijcTnG4H2NWAZuIlMbOyskbF+/4+MrpdZGUWZRSAFf8fOJ6ysv/k3MyOHid24vi9Ggs3++e
5F16j7gPXETzIk5ZPimfsn4GNHyncYszgVVUG6ioykwKlvqKnqGt3wXBwLbjt9OVMS0Z53ZlFRUG
msmyh+P3AxE0i6/7sKjN9UKAl2UIBbqyo8BKC+uo/D186uNN6dVLiOhlc+LxKBpa+zkl+jEDgIG+
I5TomAbpFj2GfDDst8qzQ4ynnju6Ji+cLZIyUFofKOlKxQ2G1c4SupEOnvzyR7fOZE+QFEfSjC20
vaIh9+zWmQXysRCxXOXqBqEoRiVq49yungW1nBx+MlehFocAyI9sxrMh1e951cEczbPTU/eV9s4P
GmUU77zR1LnNiAZuNfWltAn4fFdipnWV2RV1jsJBQizjC1P7mS1SUzhzTtMtZOk/sopT7/LxtQg/
lMGTCKcp3+azZp4qktGm/m2xe3alYjPOT+MUquDMVJg/Vdzv4IXE23iDzfXwWiLg0b5IzMzS7eXE
hrTOEK40+RZ+GkMuXtNv1hywDY+wm7ny31J1wvLCZm8BcYdBK9E8fP51RarHLoYL6gKs+zSrAk8I
4WBqVJVrRK85cH/lZUpRjkVnJ8MXvO9N/fqD6ARGMCGyFEuwg42O6y5vVJE7FvZOX1IvnhyPCuKN
lJC+E7Kop/2XxtKwKblq9R5lbYulgxsqUG4ls9Q1eOhb6CNySlofunLLm5/pP9JuL/9Uf7oKQe/J
vIOvxSY9BXcPEr9WDBpLpgk1yAyfAuMV92IY4B5aYWA+8ldiQbIRCkSSlRgZuxfcGrSAjNWobHse
h5g711fwR2tO8n1nfA3/t0PQU+qaNj8v0LAB1bVtJd76n0cmF9HEiA6sjrACjZC1fHp9aI4/nwei
gDXPyq3cgVP2bnKDsg9pbPc/ME/tJiYtpSj28AyX6Nr6fjgbjnn8SHjl+5PuxSfK6Vs/92M/AP3K
MMKJ9o7fwGwQLzPZT8khZgvtCJJY6ozEUTrppGhUFJZXULrMAtBQkQCjMpctCBJKc9O3ClF/bh3j
iDS36RcMl/3jdgX7L8cAVRYCIMSwfE+YLbR1rfUdYyt2qga4BLP7hR+Md7SOmnRP22kaeIbf6MF/
vP+7UYwckKOnFPsZNwX4ws6CN0uW6RwK/aiaZHvqJOTD40nmoU591J95ZyZAUFBEtfKqDlPR4MeJ
cI1JPquoW9v1+Ta9v43VY8tKlKJ4cLOgyYR8NBEQg1ZiIkugSu046kxTNsFd+MD9TlbLm8ea7JN3
CunwxQ5B/RZAbCVR4Hb2WR2RsLIoYftrU7uVvtXLLOtwCWIoErdN/LE7r3eeyWhDyG0TkrR3C5+T
933oqCUWlAVuTw1f2J7VegOMdBDIncQ0dYWH5Lcw9zgvuSonLOQsK3O5jeHDKRahuasuhN4QAoL9
zy9g5eXCINU+Phc2ThcqjvIykASuwvCKTmDWRtGBbGSkiIrOJA+5oN0SEtOv40Hohe9OyYb5DeUk
kubmXusMOilnF5gVfduJ6fegRBBFuJHufxl6fBLNRVvRJFWNxeEdRF/6hW242RJOUf4dGNOtQAGA
AoI7VnarCldjCI6548Vo2HEE7bYBo01WxQXJ4zi6vJXjL2StSB8HaXgxaydV3M0SkwMC5LXlXSLV
5o0woBBwYxmlwWTj147VnsrSY3sahS9mOdVSw59V1tBPR2i3GCPY+wbD+Q4YNASDkOM23x+H+Vhp
6FkV5PI5bV8XRL7mc3rGNge+MOKTKC/CznV/qexICfIClCUH6/RYmxHdi/iIFXvCMABSTYIuxJYE
We8HmwKCuTsnXVK8/BLjrZdcGMHGDs4tMqVUPeD0I+1k8os4n5oWgdPr8i2SkfqGvU26PWu6PsW8
EdRU5EBV9rSF2G1fc3Ppcc08P6yhbi+kNEgboXEVu/yI6/dnB0HVmFUXsSyfrij6MIB/2O47Po7I
N44Ux9owhHJ7BXFxj5EdpKPimWMK1hRIjPR5uDPH19fSIa5xpD7XbPUbQo8K9i/K0YMZN5+tbWYY
oAz0B5r8Fa/wj+yQjVsB/XO4WaO6Ox+pBQkGA1osfDQp8+gP4wk2rI4zeaPs7r3cyuee7rOXNmpp
u2mAqktn5OX6ywflbaFzMvIp3o/lV93tTpELc8hVe/hSpE4yDrn67f/YQ4G4QqfYTbtFIy5d2lW9
CKxqju5ruHU5cb9JNIak+0nb55r6N93Js1S99Kej8CU4ZkqWkDIXnj+I1vhGWbCAEwCBCyGhAAt7
xypN4/bZVvRpFu5/vQSmZ1us+07m518MadTtr4NS2ylrllWea+L98O06O3OQe7hFWoCnMoeFf9rs
xO9cI7NmBqlJD6qM1kR7pkg8U8LsApSNytdxMqByV6AFgN8vkPfdAtuJCAFHOQ1BnPLU5xbWHp74
SBQcg11EhlA2kcDbJ7z3EHORurXCNOmNiy4ctErB3z1KpxMfhVuIRxAR3leFGEnPe4oP/cqhPdh1
L8TpcusOtav4alG2KtyItXW+8WTe6Wo1BrUF35SQdYh5gdMKB/1CS4W9FNJPTRXKoWFaOuCF3uwj
tRMeaqqInnZe8zcYymn6f6QsFiaMLS7FkejACxv7pVYG4ciii1o7coGE9X2XGcoxWD7NbiaHTrwm
+vFxlRFbdr2wzO8MXCrbiQqG21HbRtUTeS4OeNlRTwFnvSEZW5e0OJZP1kFhxuTabRf/sJNEEBP5
ADCSvKy6jf+fRwS2uY2LlWVCjx3baHaSlpGIZaj0px7jfQN11/05Y2IbXthLoLNS9VDsQ9zqssK+
UZCVruHc+NEVaBJeJzAdvHqU7cpaGCcbBLyQxwsP2oE+isxnFCTBORiGd19TVJli/cld4Ls3kINH
TIyBG05rf7qGpU8XPj/SvqsCr0yNtnSdv6eyKwkZghA/VlM9HrHvEvrC3eJ1ZQARfARQtWxsoSv1
9Gp8z5SZWFJL/vmq+yuu2xlDuDFTWbqrJrrrvNGBPd98pa7tC31OHQl+234pmqGM68ugyRddg2X+
RHEsEtcnbqkY7n2yLBMc3GJR+P1XMZmPZIEh5u9MB8nzq14X79pIBOqgrX2iAkhleNU8FXQ9EtH0
YZrv5T1QgPskF8Sj83tfZvHYC7UhmwFo5RUiidZMO1mhuH6Bo80gc1laiGDQBP64GyUmuZo7mEIF
ZnaC5Wdig97GXB57Qn8zrDcL4KBLVSwL/xvV1oUGyCG+2s250Qubx5TeTcSw2wap8si2MRiTbcbo
cYPCq7TqevYt4SMRt2pySUqhmW+S6xzXJKXVfGyNj/TPsU6buTHquXgbxxfWr6hukQhNv3yygPXe
EaQw/ICxAEswYiRR2mewP78RrL8n/vZ1MY/uOfi3By7iIq7hb0xS7V5VllGtDoOtZRi1N8xXZDjg
8Z0igbrFvBh7e28JteWT8ZhPwugqEG15J6PB9vf5yBvxAXiRyIFkGJFaGcFvtDCB7IXl5nvrNDao
AA3qWRhQomt5xH6OnLTNxShSiMA7CZa8hfu6a3kMAAtQGkgxL+Wp1aGH2nK3XfnASePxnZLJePuw
LVGDLfddUxcwF18yS2YRYwIOMU/dV22utCwbWjCgL5zb3DwU/n49cjvMFg4tyGlJTXOd9p+mIY1c
hhtetW4ZXuJ1FNGpLksDeA3jFU43VQ3QjMlDZA/OtNmqt6/vMtBeuEWyphbiExXnwuZQH4iIhqdu
8zWRIrFqP98+86MqAKVG+/DfpQ10J1SIsx1Q4A3idrcgr/yXBrhYLV5VghghSsqnuUWpHwbql6z7
pFxKE/8owwgMep4+yQ0iI7Fe85UcB4CZckMmMPAfQEW3yU0xo16O7R8AZHcPAOCTeyqD9M7mbIW4
57++oBKEi55fO0b9YwM5MhoPr4TDonqwm1dnxQsu2EPIAzX0WQ36owJwpSFgidFcUjqLXs/OH3F9
JACuX2sr0x6oEb5N9dO+2YtRmpvfsRkGZYjbQ27drDg+WgvDqsD70ELxqFEyc7StDEmEXWpF7+BD
14Sea+WH9BKD9qr9GAIn9siwO4rZrywfJL8Qur6uQ1OdFL4BnmtHWHFrEoaSx6o/+8drlilKyQE2
GYyTaZU03BsdWAAR4rIMhh28hpX/reMPBejHGcdmSl+RQbcTsJ1WF87jWe2iVimONzHgyXLWnq4u
YV/FDktfdquikv10A60WTlRly0SP4Sy1z1dFEYom8Xf7JpoPtNSmx+D+DJffOPAL2ql9sHeC0fEt
WIJD5R2XlXr3nN9crEFY3BGGoCHaL0+Vu8ERr+d+sOvTwFsAYGmZVpsCOjXDJgIFI7A72G+xS7N3
+GdyI5KvTGo9dl9cNrj+N8yJFfkzg0/7/1uomzlVx8Vw9UeLwSXcodooqnnsQD5ZyAzSfPF6B7th
M8z4hOeleF2MSR2ZRJ3AZbEubJbROjcU0RMdEwy3QfuRWVeuW+HH5qc7ZjpW7n1MlKLSWr4X2fAc
B3GqP5Ufm+wl5r1Diri88DDFOyvylwftW/zQeP1PVHMp62aQVQX5rxC6TCls+9B1AkqwLus6H1jv
b640fftQk4mpm0gfbgB2V3FACHudTVX5ysXC5TYpT01gynsKE4eWpA/ZnTXW4MXp9jlePANJqN/P
HR4G3sbg6teFC7LGums1Yi2HJrIsD2nxGE3kJTFHEc2UH28Y6AdafIwJpZLVNYx0I/roxjHtJCjC
9avUIgmjcRi9KqH6Ypua5i4tE4IEmT6995BoMBDf+uLAIET0z2AQEygT29YYOeC6BUm0qKFmkPoM
7eH77+D5AVf3e1NlNkB6gvPPIJIx6GOpxjQvivLL+397DRaODH/Xe+u2rspG2wpet8w+z0Qwt4+g
s3dpUgZg4OwSsVwQEcLpsmW3cHmdSvP47X2tjyv+olAur5tQnfDPoFuqOMOpXvWVUixDqpYhvUjP
l8bQSbTEvdJN2oqSVihD1CL7sAiA0RvIM7SQ5lQ+uGZF6zta3M58aAM2ZhZiyaF+CfWg3fVgMcFd
mcKHVvFV8dfgMPU8KZL+3G+umvqb7MdBKs5DKkp0b3csAZoe4ooGycW/km6erhqFLxxWRoH27M+q
I/YZzPvUyacDXkO+fjMCdk9vwPgnz9cK+nIXZ4sczu1gZvyx83EakTS02d+yIOQRCHKg2tLI//Bn
r0T62LausOkqYiQR3Hs0xR+3wKTsVMsw9wOwy5jnv5It974quD4npXGZ40935Q/6lnkY/BTUEFAw
BpBOw6m0/JPMguZYKqB90ChD0trg/w3AyNxMDaEQP7olZRBMI1JWcyopAXNF/KlgQ3sYFqLg9cnr
dmilLHPb9nB8ZmRDyuhlfGnr8jBA163enrRxVA7Ak87bBStffg8vkJqusltyHawqckUKMAlslxjm
OVp1Yhj3WvO8O8e4PDlOz838xlgVppf3XteFx32+6REil0aJH8wc2q2p3RNH3OhFZ20PQ8nTT+jm
AC65myIwhQhspFT8nHpkqtALyfU0XYXGPolhfxFqS6ufjj66N8+PoypJyMECsyDP4iQEqvY242IF
NUx7oV5eg1CAtWq5P+V2t3cxW9Lu1qs41P7mS/Wu3THWdO1qKsbpN1te+mOprCXP78lcuEiKE7b/
FY9t8EC3X4d6WZcYvNX7QYWV+fc4UBPcq1fRHf/Wq62zlHRoL2PjE6hB0pXjqRDVlQ1RezL0lzDr
Mt1XML0dXaPEOJq8oYKPiODEVrlyHu5uHzQxlWLO/4bIHWSsL4CjXxl776fatWCSLKH7/Itdg6o4
JmBiEvB2AtVfUmFUHfLEzw7YPVgInjjXWFo4z6wL2VhypvyXNnWMAWMBe/bFMD/Ee4uquMgloY/C
jk5XE0NRyj9zzy06G8wvYrZAUVC/L18Jj3QZMJvV3bjU8KJW84i0I3Eyu5k3KvJfaA97vOm4XOXl
Cn/WcHJ0rSFA8dhni1nXBKGVlpEuxtSlOkeL1jnGoJUtWUe6D8wUFfEFkXBQOR0dfOdXqS/GfPux
lnVF279UEAtMmDBa9FaU4gWXrGZ2ACPfHnqLkbJHtGkFlqg8sGuWL7BaC9kj9lw+mYxwG99uIEQD
nZ8ddUsYbyDbVjGJGpnjp79WiiXv6jldHg5L+uyFw2XehH3J4JznmB4D5Xk+O7C4l95K60jJLsoL
1Wx/xPmRelTJYDn8ATzW98vXoydvwIgm6A83M+kIfwINhHV9W3wlvnc1RpVBeAbd1GqAv0Q9+Bnu
JahERxVehApPvYuMDKNr/aFDiKKXJ3ncImACSp4w8ZY/rbcPcMSFc9SlYpGJBSKlEN5L52CVgRx7
80ZaabJx51Doj4dYeFHrzGzZJAsx8aq6sBXJk65nYbs+xEHqgdAFvB6PEjrcHXG0l0O0dZhyRO05
Lf5cca0t6kruga/vxI8CoZ5JTjtq/j70JvUqyZ+0BYEjVnmJdBhYaA4sJM8mb7tm0DXQJzvGX2iE
4uUnW+evJnY8j6YAt167nXsJONkRLmzYPUXXT8VHZ+buM4obU6ksa9gLw9Ns55hZLo09Pi4ovIIj
XmUAMsBBNqo+eL5t+yi/1AiVb4lbVhZhgrMZcrASq3MvSYlnr5cFQb+nvMiXE+PbZPAWZqFuqIFu
RiRSFAwOCGN9MAaSkEiHSZLb8AOGvVKO4aokbO9b/wD+3STdNx8sf1U5msVBd1G5NI3dm/VBw5HL
ar/dsRmzjYU0xQOcbNBCcpJIHO+oZ6TPnKOkg5AsLuQZvysW4D39ryLAcdS/8fKXagdYkyumgaRF
PExbnX9kTicVa8maLb/l/DwpS7dBtOp2RnXSu0TYhL/oS6nC7GM8s4LP4on/hmfij0Qf8r1zIAbm
G9baLK19e/PT1x9LFHo2GR5Yll0lTr3eqUiJX8kXmwXUCCKWUOxMNEpoAw/fBoGA/fu+OA2j3Zrr
6lUgk4VnJ4i/SG//ZfIWhSsxPQLJ4ljJimcyb6bv9NIOTyg8VKXjiQvS+SnhJmWyx8NPRQfD/GDO
uqYlZt5Jk1vuSllMsh/WPSe6rasAk3D1qMQloaPAy9iecLtKpReCR+UNLChf3Kq9epwBrUO0uaQ8
loAaMYIXZy4sxrsnJGE1MWQNWEvNJ2+L5tqAo4sqK5jTOQW/S8WxA5NQ2Q+0DjlI1xrbTbVFGKQ3
rdUOsxBEa0eHlcYRJ//cYlrvJkJkLlW6bwsSN5EZb9mjMqpycp2C9FTlci24QyXVcvkucGKJDSkG
Y60O4+Om4mP5iBriQHRWu2GD0d/GEqI6nmwMWdihPlBQ2HwB7OfiItJ7YKUD28/+4MnmzKVKF2Dd
DhI2L0Qusmhv1Y1uanbU2r6qATKD4SjVwFVrHyO1lLzM48pT14tNKPbYAju29BFP5OBF4+pqlmks
EyUGE3xIV8GI2Fj2MPDbKVb7cftJd1iTUuEFAoTvA3ZGvLzePber6Vwn3NWXGbZiwc9tREbzvlgd
skhd8LARHujPdT6xmacOIIC3NG4OjbfPHeFK5Zt789Jr/j/P9TPWU+AJxtXhS67E9IH4BNm1qeBN
Bzzugb3RV5koepkoyrPtuNmHPVmvwUpMLktyruug9rK7DO9jMwI5MGRTRI+2LptyvR6YIkKOyDg9
FB6VmG6sNfn8TnGiY9gbX5gDUBznGpiXFqzn7oqXEVPTJtVB3s/o+LkiDkXZcaLrqPjS0tcIzlea
WcRxdcqI7n12B6wF1pPiiSB+3HlPhOSt6cP0Eb2d9+X1hO7laXSD0gZdUehg4Cd6gAelewnEXAsa
hipqHOf/XBfRneY2OzRyUq6oDJtsttSkxwK3f/PjJqxhXISzW2GY+trtW2vMknzxJoS9L0k3o6LP
9QwZRtCDxlIn4hFUZZ/nvqiFG6EaonRux2gZNY6OmF3/hWlXYpeCZiZ8zg9O8o/5sNOi+aO7+0+t
jhCE93DirQuQ0jVqEakSnPKp3JjH6DAGvZjv8nTYRVDC+c3DsFBmwj/dJSwagAhMy8ZMwKQa/iDt
ofqZJ/NXdwLN5PFURoeMIuIHYaEFTusPENgndp+JxRWq3cd107RoOh7IL1BXpu9GQgUK/16MzdbD
iM7yTQrM9BMv/N+VZ+jzhBs8P2Ervz+GoZqpInsATI9oxqTuM2ftYsqOABpKIXKRKEGuX0vsS47C
sAYEb5HTLTwuchoNvf9k14WJP1XWdKmyfVD2Q1HBVnBwiKszWRcZvWKg+hCFHYmYvsNLpxrD++WF
yXl8nAYJfZ0in/SfUGyGn6/Ggox/MEiE23lPHQT+3neiHo5W7HVyvaYHJqRG1uAD2lBM3gHvhNuo
ykd/WWnaZevfSFjy/sv4Y0caHldeGBruM3WineYfua0OT9weagmFlkEgAOBWbW9PPUNmnr7zReXi
5BcmUD7MFyXfxL9Xx2u09oidS8S0EHf/cvxYjmJ3x1S4pQ14paXms7kuBTx75zYQ9zAAYrp/pYRU
pdy15oQFuD29vQNC+Y3QdCmleIUepZ3se9Cop/leNar4o5ySqGeyU0YjZ4l1iic/qOyO33NId0EK
PxkAzIst5pGglnCEhacZU4uyNCj6Q6GDJbN6JYTjxQYK9Xcec7d2Z+oFvEnA8fnVFICFBW6XTIPN
K5VONOMfk2aXQuAfr6QUEQpOYI6gi/aEXpu/CPz2Bscx07r1l6F94gBHfUdZoaLqqQapngff03Wo
yVzitbdUmfLihps6eHjlPf27VC+ilUUjmeNizqnm0Z/i8VhRMDRwUvYQ19na9MTA24BUYZUm1Ysi
1bFrN+IUmFk3aD13M04zVo6UJ9kQEemOZ7h/WpAjGhJjZnu9lCMfgPGmkbMfaImkr6DvprI3nJeO
ZsyvtLFDdayRMEzBFzPNTN6uf7v/DEhlnCI3ENNglOgmUpHm1Vsvx5hNTE5U3aNimEbmt8G39eWm
fzh1VmoeuFhzMkAWNAp/j5T4HaHUWn9FYHsgqj7VKpU4FV028Vy8xATV1EcBpJ9ia8v8MU6miOcT
vYd9G0ITOB627nnQFtbZ8P9Kz+KSk/SWDO32vYcqBO/5rwXijiajB2DV82qc7pRpPCZxMCapxZ45
TwttYKcITJri0c4WvJJMAWQBhC96sbhAznHgJNoxOFv/pAhwzkVkn+Fk1kScEjDNlcXhppfsXCBs
43I68NaIu+vHzJZi3/eTEDndQ/UrLQHkBGBxKTDrQjuXJ1tPuWk3QQ1NuroUsHUxpg+7gQ5aDFaa
YIjfWvQgxMorQwF6MxZ8oB/W1xVD5gc0Kl1YvGYc6ebwMfeRmJlNAbzuISXYtZYOVn/ot/I6Wwrg
e36jsqwirUSjEVeu/gzBZRIYqAUmim2K4L99/gnE9XTWTfwYuJBjGBYVt9kH6x64OR3I3dwC/hJB
aFDTSHV3pI1wD/d3xIxWEpyRVmZWSf1cYY8Z4fOvjnFjmx4GADu+hDQkxAQGbAVcA7cSLqmLvU5j
tVDMJeTSPlz0yivq2UmlHbku3l6WDs+CRmSma1/sYIv3WVZsgJDHgpjdbvArgiNPQNptKJ6qUeRq
ZtWL/CdEYl3CyVRD0bKXpldyVYWX5AcecoXgOY+5HWpwka7dh9Rk8YfvSMEd144mM5Tcj1Wa7p7M
LJ3lTOzb0dabiIZO0tU4j87zv57o+MXpWq+aPP1O3taYLFXvORxFt+p2iAeikS2wiKE/vwriW8r/
fC9wlwsBhCz7NAuQpKqLLLEqihx4Np6TwSi5wFo4oPEbklic4DULYWzGvqbUrpQks5Ql9CL/rihf
gffVqJM7OhLsXhVi7WM+PnvSEAxmFBnVqYVVHe/g1ZAOTb9LQFyYCfceOEkAUjA8Z70kdN1AD1Tj
L54+gnoJCtnzsbLlKc00DmK+8Rbg1ch+yJx//pgewdZ4oC4xRH7XSC9Uuduwbn1NmZ/VwAiOBTEY
fwX/AkIk32W9oNDwlhoN/43117FfUBmtsPsZF18Akic2+9ItbFJ4FdloRjCae3wBWRonA+9wekLd
CMl44B4eJunB6cJMXzq+1ItYMXWaw70Z4XxFd/GbxhfD0eDLbgTKBLkpAbwH7sYXMoQyE9Tj2ybC
fMMwZDX2AeVHSULkmIhIGHYw0+j6c4Lk2xXXxaXYJMUhgNzJ+5qnJOYVlJ0eD09/ilMUCRtJQrk6
mhsa2ExqZ8i3dqXKfgm+8EYDjnRtHmec4ExP6RJsyQ3Astdj3ICbI6t2XGTi3N0A4BUgLmTQolXk
DdDBMRLN1Carv9aqAFtV2e9iV9g8vxSbzFpMMS6e3nh/cLXWeSibCC5u3IjFz0+IMIBAl4E2bs8i
rYwbPFpYweZyXNInR2jK6fiZuCTTNoYunHR/UbXqllZ8KoFu5uAU11UXKTvz2XKkveGEl0Ua0MYb
YmfEBkzbp+rmdOOE3rCD6cRN6738Koi1NpY2jrn64rzG2W1wi7sgitdO1db62d77Lj3g6jEcFQVi
/VL9PRAf2CZBDIxBrk0GyL4MAx6ARiEmU41susE8V83wjww+wCMOgr4HcYo9kKODNs8G7zD2VHv5
5nDmIc7ukG+KUN9JuuxpxEY6ewrf2ar8MQIBx6MeVGseWyYWQqmZB8lCGLKN67DIcMtryl0Daskc
g0CEBS5s77WExQRSw5eFQWhGXkdfapDbaCTpDPkJqeDbgfBX8cfKlzjhhBm94+HEI4KMaIXFr2A1
SN/SDwJBtLHDYj+DZt0SLCNvojGO9DL3b6QGpHyyyi+GyxgTxTTw+2dX2cT8QdUenQzHk1kx8tq8
frDL70F58MDv1F1iiFbZpE0fsH36gjwi/NDoEi34qq7NC93FV4CQCmJFEWaC5tf4Q579CHyvf/iZ
z/tJIJ4eHM4TuIUvpgKe37ecs68R4PP2ePI9/Jf2a6hkvMHHi7m3WI+ajAtXFi9rQoS/T9jHq1D9
LnlUYnrnHKo5c+qiiRp17+oblpb4m4of7YabkvBulN85RrUTHsfy2rBABA0FbxUfZ/PMP+nR+igf
8iQChtq3TvB4EHB8czq7SEcu0v28ruqEraRJQCV042JjG6mrE+5FqjG3rMjGWFuiwUP/DrhFshTq
OysrmljCJDnPlb1+Sc7knY8QChE9Zlqqx0XpjntXtYPHsBUNaxvuNuYV5YbfS0xwreYsgSBhWG0h
E4D+adocl0h9UownQT+EAOhCKx4wAkMt8y56eUviTTKsmI4jwgOP3kLFpKzviYh3gyN3NENWOKn0
0sLR0P7OCy/L98Ty7rse8KMluzH/hs+lfUAfkihCUe0zn/oFBdr6vaEpUcTPVUwcwu6IzMF9nrQY
Fi1Kn//Yc1H7b+3RAQ1qvrjG1Xvnubg5s8TSEUNzDKJkqUaNyeKrtFf8Ema/6l6bxMk/4ShXbc/b
72R799X0ry5f6DapzjV6RBJwptxGFNJQ60JhT02BmnaCJKMl9x+CkBUpPAUoJBy0amJAkWrNw7lE
EDmSZV1R7pR1UoTomJa/brVjNhZqvzRyvCwpC5w4V2QRmpaL3lPWnsN0CMQ9eqMceZz0wMMuw9Ze
f4mnfNl1kkBVvf3QxIQsLLROZo7l+osTNn93SNcHgVxPbNESIrRz5DjEGBaFSvAPLi3//K4XzDU+
hIg/UtFUcwa30ywLGrDP7qQJvWcpJFdJU/L475D/iQy9gLP9/VYoN7VEhtDQKjdfQX0b8hNosCuM
T7F+v/nUoDjoo3rSG+K4oXVXg2LaDAo3xIE1pKih82PNRvC+AJneQ26hMSqDgtxiedK+dzCIqz3/
4T/1Vp/dRuCNwbEhutF0esjWuTp9ESpY5C47vZsJNFCw55ZrtWZWFHL1+jXqcvgTGscJbLiUr3uB
hzLYJn0zkC71I+a+Coc6gqEzjrPdAjhoKT9Gqv1cm0sjV6yF6TQwk0qyGjyIxc1luHdqrE/3CkNv
L7rlqMaOQvDnC4qhL8zEDsSisr75jgL3OYOBFTpnbB+1WgPVTZrfRp7lJ7VyOhTryf7RMgWh0WUS
p0WYRLSHUcWSY/6bCJM2Vq8hR0FtJuZuRZugBCESp5ychio5lKFmg71ykmCYzUuSnib8eIXfUQKT
Z7HVuPXMv5meaJfVaTWABTTbCmnaXSVqpMf15qL7W5tv7rFV8VZsq4UWhILRRfDba1tn+7RIuLYX
fB6MF4Z/5dm/lN6xAsofzvKLWuLZs8dN2nwvSg/HQ/O7JJd39u+dx2V855+pqGO57QuCW6PaMzRH
c026ADY7Y9gu1mjkcnbxjNU5EjKmVjY0KPsEidvx4jve+Y1V7IgLH5pPcP7++50sosapcKOXuq/y
u4cUsgYnZLlqHlDXZi68q3+0pjhd22PF7NGghxldacMdsnwCwciujNmwAMh2Aa7g9kQwMVo41eL9
y2EqA1fdaIRxxlRXMgdp1TNgjKkELgxmFRxoKV+uI1EmzlCccRiYgpt7T7JM0TTYPuetUMrqii/J
AyKrU/rfzzAWnlQio8FR7vZmrYP2o7pP/ON6u57RfENqsdLRmR5cvgbWT5FZ8/cbpSgH6PqBf1+x
+AlaoGWr3tLXJHB0kFxHPp5AtXvBluf+fuVveLZCzTiwIRpU8mVQsnZIKRR1vvPf+dm7O0OERIzb
GVCk2u/5+TD80hTujlaJ2wOMx0yCv+1sdXyvHMAAnCudhdfX+Sqbjbg/8VTJRY4YGM/UFTzlpVFI
x2tAola7YuusLTgSzNTAGy0xhHkjthYUDw9hXAS9YL1qYR3cvL8S1kBmpjUiGglbw9qoU/lMRWgP
c13oR5mJYGHUiD4acDDm4aBrLCKvus1HiLcrzaIJ/7cKfwzv1480IjdwEHFZQd6MIvMqED+Syi5Z
jaKHZxQEYNpPNZfB0kCbQmetfi5fnyi5OjR40hBmZuzPLdI4kCAflOmyOGs+bs7sUwMmVAB3GW2S
n3Ge8teMfaJ1mSWjAhI6skoKxkaWOitbUwR37InhId170ahOEkXmk4DHubr+VLFn1Yjgpeusi3Wt
oeFNBvbJQ94cVgJHNLDWARCb1FMvvVZPYLnMoDaSFxpdWJjr17tAXX9ZBY/1zI+hH3+RkLup7nVn
FLCby0n1v+8xnKObFxJknissTmXLllRNHMHlhkHphgNa+25e5P7Rfaf3Q9xwapxpqTxXHO433G+N
bUJqb6iCXCcuDrhIiRb40valBqSy0Xg84xO4WNBHNenFsq7VAPZnmYFb3cIAouKb6VQtA9w2qWwW
cxdZB2Fkhy/rbSo0sQzLegnhJ7qkUJiqLEVdzbD3mQ0MFzs9S1TcLEqv4Pjpa6AktVGWqu2qD+om
TeYFoLo+ZMWpYYoUu318LsE2kPX+w+REvoiG+zHy2Md8gpd2vpDpvT/Rw/bDmyn1CqRr9koLhX5+
pzJE1W635goaM/UKAS/h+Y7bbIZF1UDdm+tsutMGPi3suV2lNIxEssCKrtt0apIbnCGP4qoafCLk
3wOyUiAUqJjrCxSpdkk1n2O4Ij4QMHdCpmyD62daNSEk2q+xaLvvMZlWYP6L2tXaMCNcXu5XA241
9l9gY4fPZeD46bLIewM7VoGOfnbLsM5b5D4MS66NODmRUT5QyMsMG5Memnv3XcgW3f2KsGH0aoq1
qxXPMKDSH6zjzvnJ23iJAu/VUMzEn6osPPwv8McP2edeuy3fxWdf13UYV818j65qnVTc6GvmlIeF
JJzPWDgE7FeLLUZhn53KvvRLwizBL5UUwjZ/BAz6iqWmoLOjKOZH7E8X6jzBbHkju1VmmnuqqwXT
mu36QgU1XkKQr9IBfnC+/W1+2L4kBjM2dQJcsrcEZECH3MK/gkg3uFZsbP4tsHuKyIRpNiDZ3xxD
TicGjhcDHfHGqkNoYdWNXfGqJ9ZmXDa/0nGHJ/yqRCQAr+9a+y9/prsqTHtjdB0lUKl4fdJ5PTfN
YQx7Wge912UKWVVAiwvoITGwPz3J+r7vkx6X4Qh9oUARyW31pAWKBYMvKCAQjcW8xn84sBYKM/Gn
5PUXBaduLjueupq+oB8la0WlN7t+9hLM5cLUPURyvRuzuK6GpEgUB9V2HB1MggUZuX/lMcuF40I+
cVVSDv3feLrY5BtL0180tifLfFd7m+PhnV3Lm3BR6SGt2i6tz7VGKV2aQFjkqiKHc6bhoI+Sql19
7B0QrU+BaADpUFUwkTt9EmSvzDZKG0Hy4tku+KvYkZTctypTjNbEiIAztjXHsgr4Nl7vWrdOC1cM
CO592IqmyDE4haRs91+WeZUSupuGBEcuHCyCKGXewOtTRlSbvg4ZRkQEe4iO8mrFDdXYpm8Gldph
5OhmifkXMngIvuKIHWtEdx6EPJnAVvRZRaibVj8dagKRPL0H1xVu9MBnAo854URVXrQ9tjFfrrCG
0FGsL4PlGqumAD3ZGEJAxxQT+aBJwdzk0/8VuTF80U+zHrk1M+FURDmHqKNVmG8W17oxOY/1y6Ip
ZYmqK5ly8m2YvpCukDe8QUwxLRdsKFVSPt9wv5lEu6XaQwnn10DnY5x0vOGwtoKN8SVmyDQo6MBn
PlGZDZRtwdb/blOraZSmmkl4MgwAgIRFy59BiOvRDbz/dpdU8hfTDkMf6Ef6OiEvP6dU0g2EXtBI
vlJmbJxSAgvR+krJ/cOhimKdF6QwIwvM+8jx50F/66q7HVmiVZ5wfma3soExVtRfu0KKt2q5Vn7X
gvfaR+yXxw/2DoEJsG5mWT1+u160rWEHeaNUtlteZNn4m0b3whh4225v/WfKm2TVnJiTYVzniOSc
DYzg6SPQSh8xELBalJ9mvRe7RZEsXpasufj9XbPxdHmy7yoQinBOVPaAFnD7LPAPy5sQesM1/XcJ
CIa4CiJF+PzJ1Ybtj8FMFK4IQ70nCowjVnAUed97wtYHZs/eoFITMQE5gJ9H8u3S4TwuS0IrfJCe
EXFkS/20S3W7PZuCqTAEw+o4kjhDX6XKcBY0EUx8uDDobrtOGNFnXASIA+uKy+mJqLhwRMDGFnr2
xZKMEC0qdWjYpXSTDaht84O5HTtVLRZKeGO1ehYPs4lfoALhWRcOXIB+I7AiwDIYvD16J5tV4+K+
YsHrcR7HjfAj+FBrwv9G5Ym/LN0OPTukYGcEfB//MIOu06wTdf4VZ64pHRPYOo9cM9BxjaK+oBh8
pQLVRINavYmcnDuE2pAQp0VrRAWmjpFWy1ef0jEtBHZCAFeR+5F2T7zwRYpmjVXq51Bqxx/+cq+V
nROzdmBLhySpW9qwykW5clhAM2HrP7cNt6RdNfAqeZEb6k9OZFO0xyCe5uAx3mcs4FFM/qZu0oHC
U6EuhXjwyyyMyqJCHmjdtH1bLSlLpNZhoPfQDhkZUYe/hE4c+vY+eyzHCf+cmTuBk9gO41EeYUn3
FB3UttF+fEM4TtwAXDc9r/rJOBjC7Keg0QArtuUOJcT4yn/ydA2YEnK7rzt4NMfTWVR3bjhg535i
ltnTq/MIPoC2eIcuwLeOff8SETB5pPJJ7QkKZct1ysGmusH6VM30zHFW9uWqxMbOrqPPSzWnqcAu
0WTuJCrBrsqk3q9y8o1OWfq16VzhUU7MSbWSvj4ckCc+nDV16P/QDJDz/Qou32/wQJG/hdBDKf48
osT8jQjyMflP5WNVobRK26v01oRLd6FyUkkWNJB8zeW3vLFH1LB2Ar8zUUq7JnVJAkxx6io5UTVO
mFPm5F0SutAHZaB/JyYMa/hjccMmRaqgTxhxBBSSECr7XZWSDkjVhYTDnRlo2eUBA1exdZs/sXIM
Z2aTXTlLeEoSJb7G/1uB6qKKwTDZW0sJbYFMhxexrjP00a4lnrLe+5AzUtMwFzqyGFaFnkeRtbsd
UWK0DXsXle8PioNUxmlqUwnJJ4bDukUwd2UF0BmoGAfWr28uY7oA+xMaBfGi8fjtTTr7GP+V/Y5q
1+sYm3o9DBH+ARzTnNWrfgbl0G7W4VejDEDXp3T+gvziaS7Vi2rLV3MmGlodNP6xLB7wrJeiXhcp
swq9zVtJ6t2G6xyTULltvgaFwFAXXg3UNiWxTEYdBNVEFhq7gthPQR/GvnzRYkhpeBvx0Y8qZ/1X
BbW91W77TLmWbO247mO9IfPFJktZreIyNaUsUqqcqZMGkVq+xFbzHOc3QVj5RvgKv6QqiD/cCCuk
sI4KAQ8af2N5m4pK04uknRXfyT5dsym4WeUecRWAQftNOAWtfPw+/Aw1y9a+8a/gQXMwWn0NFmpU
hLtj5tgmtKiFB1TTYsUEUdDZKYgFcE+HsuEyrkoVSRKkwBRQgV3f/6UH5I9DClX7N04Q92VG1r9s
Sf5Km7FvrrE6OcydBZsGUmBYkgUzXj3MSur9r4DvTSQR3IbdJHJ2yMB3+sE0kTxCbnoaS6xvFQzy
09+4QTwM7kIk05peabxzaq1e2g+hMDUBrvKKgdNb67HZEM/9HiX28l3/YJLMPldksEhVHe3aasdF
1hS8R4MxsR8+iswQkZwasb81Yhrm2yHboRsaXHgpKy3h5LXOK8SyQDpbcQxBJqG6RWvC8TB7QS+R
XF34EeQ3OHBeNVPfH0iX88FTavmAntXQyx9mcEZsSOODWRLgRDONqb9OfibUpQQJrvto5JPkXCuy
t3x2LeDp/Ee7LWJK4AF1YBfrn3RAdXKsHrqcTziuSapuEDgUjMF71ai53Uk1V7Kz2x7VQhuAJ+bs
8b8b0Bo/4RpG3lAoc9VeSQn9y60+R77nS51X+YXs1t4aO49PrjJyyRYcBpNlZaML/A3fjXEh7lUA
WzeYaIGVMCxc2EdiuXG/qOpQR8KciSLATlkVP4+otQC15RBBEamyAPT0fGVftc1sKGLhiwZpVXgr
Rm+zcubQRPWbahD6lc0PpolXlZNQdm1VlZ31F7Jd1vkvWxx2pUYu3GUGoS+iZlEV4xGSHSJrBg5G
/KU2d3T0P0HhYu++2EVMulfxndPNlYf6WK00QMFH4znprIHnyxn74csF50C+m+MLY34GQsLitkcA
TLI+iP70+FYI9sBcH6KHIAXnoZ6UdqOm0jnSlNv3FKRZp5fojX0eVBoFbFmn/jh3aA3O1xhCEZ6A
gqLNhdnM08lF9J2nDMJdI7zGp3sb+mzk+g6iAOMT8MsyR6TK2TK9U9Kcuz+mNCc3r9g2BEnL+jDA
kA7eVS5kyNrPmCKnNH4nWXOAM/xC43edpw/A4NVuVM8l+idKeibLYcF348G/NXkpbBbp5OGb4pIn
uelOh240BpQ106fNwaRftYa21tcZQCDgjmXNvVQLfqdZRmx8KlNM/uHejgka08ryyDQnxW5sruL0
MS7YnnPqHg0oT49xW+ljY0k6eutZUE0rIzGk/HKE5lDzi+5xQVUPMmhKR3Dqz0ZL1/WlHfbtiZLg
2i8n3bR9JkGjv5RSchOUZEaFBw/dL2DFAOrQpj2vmTJcGER8zyoHVzvjme4SomkO3UF9f7jLFmlK
e8Mia6nX/b4G+ZxuIuwsodDPwsBEj/i0yY1W8QcCgXiscmh1JXFpWZpR4V9NNxO5D5pKWWVw4l8m
C3nhjFqhs1SAxn6xKdESBB65koUb8hV4S/n1I3Hd9ZcBT7aXQyBxfM9ZrE1AP/zfYEJQDcdzpGBd
R0+MQIJ3T5qe4MH2A54/ICTtPr26OiJUxMoSZbVqca5HNAomR/wphbyqMrO3Qjb+kFYpflv+EzTa
gC6+ukgWW58qJPBb6rWJMRNjRQG47TsCMnZJ3IkSm5s3Ll0CRygP3LIerTSIRCu+3/vX43YXOSSC
5m8gyVAJljYD0pXWe05Arv8b4XbTamhcmcJ0S1rDHMlgImi8ITn6ENLbbIvOK/+QTolwEstIBCuO
n0nxHw7dPflmReLRZ/oJ5rEt7PIF/3OuR293X7JLK386AULmYgd+ZthhZmKrGoTsHG5mXwn1d6U4
7s7LvRHFx22J9TsV4f7ozRUuHJsw9y/QiS4dLdacnbl/RnQ/jccGkpz2KgRIBayUF0ZZd7DyB+yu
53QUO+SBMfUkv244Pt3ojEZwDVFlOIurDSSXyXVNo3kC7uoDRPVypfAAATN5qpyduObGdpIUzOZi
HvklHYPLTmjFR5WrIVfa7zbNSs2JLK/OoiVpsJI/+p3KJYf8lyR/KDV0WzEYpPbgb/KyqcTIR+fI
hmaVneBcQ1DIJqpP70jiqVcNW//iWF3DFMwKOIIKE4b7aG20sNG6oJmwniMlTdUu5FWAH+PkNNyZ
a1dnNKs9g4I84U4N+vPLBqu0CEGiugK1fbWoGsmizyRMIw7lNyCFpPQcYGXY5+6ovMh3aXfhHOXc
9CMq9ee5vILkBEk/tshF7LaP3/sZEqN5bSyi9QhDRPTIn1xYV4uyxE0hr8G8LTBrn69w1JLZjJE1
ocp+XREhyNQ2e99bxlntwzbLVVI2rg3GLrRmLj7gQPI3wRrEl/j2n6yUfgleJ2tWUrhru0VgkxmI
7wU25Vn3XEuPRJSUdEg68VmPD3pXFFVPdWN41jAhLiX/FKBXLAbKf/Y5GdKE2obFGLbyhI63qcVb
GVrPftVwEPGj1KoWOxyStQZ4rcq4JCoCAnHQIfd6DmTtIUYAAiXFtkwTF5+p+spI3mk97wMlRCrI
qpKRXgLUBQSH7idc4U/PbwmibYgKRLhMt4GOd+cepPyOcuyHYPW+pR1RHSknBqFtjG7Y+UbG9coq
1RfsVhkhwwQvv77WjWmJ3StF2wlyt3Q00JnZhRufHThvjlKC9SlslWnH970XUmXHSYMAcKDrIwMw
7Je9YG+vSIw4DyGkqS+U1xl8Ox4pV8i2eBwiw3BM6MxKxbVGGwmcEPmwy4S3D5O6Ka5gnxdAUnw4
4MCEP2dRAJmGDVGmvU053M+X2/kFcem6OWbLvgwJIqJT4pAUQm9jnnhKg+06TkB9xZmU5vdgg4eA
UEHMSqdSi3JWiMQXE4ZJSQBrkAlaJjssEfww1EQ78K3uhlHkoqKAxvX5ZC+ok9MmsRkmwFvZHvhu
kYoGATnJIB4xZVbxlH/B4lxcJ4WnEeL3CEXqqo+DDDzeNd1TOeQjln0Pkle3Bqk40FJZoPwvwSg2
QDAR4tbxjZqWSPzZ0trnLPw6RVU8oN3ItnGX2ZMNYKK17iDrcn92mcjLgNXw0qlq5wQPrDz1YfTe
guH4ED57iIMphVkKOABIYpxJXTDBcZKNmh30eQTyEftLV06DnySSAxU2PIAuu7/qtjeOvNV+SvLF
hI0ngQjmHXtsT+PkJ8Rv0i8OiGWNMRoXnI4BORG5sHXLQZDJkancJ/t7S4aC/P8B6yUIXof8h7uB
YXyMHGtrrf2Eoe365np/BGeEocatIABtRYgD7yKVOfZCrSWfKU/XCE+aOv/oGFig2nh89NGQzi8O
kfxFSGm956oKUeH+Pudv8+mvec/81rXsvYi5dORel8HQmhlgy0mlvSzOCYQGKMMSbFbSsfiDJ7K7
Zzn8qA0KCnzdt9TluznFiyGX5K8u9veMU8/AK7oHQU2SE9OljR8pwrRvMkbep0zRHMx74OnnCELk
pYEINd/njev0CfJHfeetw+Y5KrVeBCTCfisl9OJJLY/m/+J+MoNfZmHnPznDxnJPKf9r8+a+LYd9
u6xnKgTmf+onWt+FACt+oiKLwPaNdyWPKHaXwE+qI0VAgcx/ZG6xm9yDqAn/m+pqsScaxu+pOeZP
GJ70wTL2alttZV69NQlWzIcF6psV6l/z6ak7fVraZ5ivGCJGfuFIfmgGp4YvuzxgJuJoKjbZuqsa
DFwUZHXjsJzshnEI64iVAny6Y5RWwefOs+SXSjE+mCOoJ2H8/JWzc7lXyER1eAnThopIBL6eVfmN
pEx8VSi04EBnhQdXSWQvwrqZG0/iURyRtm8kQzaLqP4RdraGspVlkOsomQAu0R1cUN80VFO8tCXn
3AD1PXQHvQOnJ00qjirqBGgeeFIN8HVy38gxMiqz6CSnADUkh/uW6zVXGTC3h7LD9ayXw0veo3gJ
LBKababXSosPAlsRK4NfC3iWOU53rJcsJtAoxsglC2k6Q8GlDrFI/Cnb8ARMsLxlcQDO9Z+GGAaf
OzTqrQ6tUpbMB0I7qAiGWUFhsT1DCTVGAKtcU5au5DS6tT/Tmy4VkTwRPeoGNjRcl4Ix1nZcGcYJ
NTh7XGm2I/A+jLI7Ax3/BdqfiwkpGA9plp28YL/TxxnG+fyk87O4wAd5FKKAY1WJlTDHP4ISKC9k
AjUYsFaB4xO1CkJjrdNLLmjb/AwesKBjYR6qxGoIK/EO6/2is2JbdoiKt+N79nEJpcXhNfnvBduQ
7EsNCHNnMA69BY+4iMEbElMEnBw7xsdoPrZBTQgTxaX+EL3iZax3vJSyVYeQRFuH+LOk5f10KuIU
tPM+lkaOgOPEf59hpCW1PNXMKA3/6Qbadxl+R7+YEa9Gs8XmpGaBfMZ6e+OKTYmKWCc5JvzkIOEX
eOf+BAf5i8QqtIiEY3TPL+HMfbcfe2Gc0L9nZQGaN07QrmBmbVhELRN5oPbmc+Y+FVJrUo+2nlmh
XmWCsYQJEjuJGHvhOUavGnxzf6kwPpqjF8u5GlHI0tbOGuiGoU8BQZtnuBgbLptxHkgRF6Z836JP
cb9aTI1dRrkBwNdfumiDugHaDtvP9D8jsFWkHMLP2Ttq6Vd2Aj2oWFpYiPPSmUOjMha2V9xLtQJJ
JNARMrI5rOmTtUGvRq4+PqnPxSA9aK3IlzimXegnK50ZjtWFekqT1rcQ/J+DTo6EJPNUo5LcS83B
YxavSmaudVeQVAiWOfl7GSGDyj0upvT+Ty+N4dCKcgTg8O8vNNKE0cBEcJstyRA2mucmXWAMQHLE
w9GVJLBbS0xyE/tTKb13Ap5eKkL4rHZH2xxHE8A37EQLrWp/fGhR7ZvljdtTl1ZHXpYK26DkXVTG
azfVEp20+bgzTYH4REQ1wGxEVYYJPOMtfCgpTNVfv2QQthbaDglKPfcoaeScXma6OdhzNGjD/Wqj
BuYOglxeYvTZUAEKn2Y3gyUdshelh+xbVVns9/YiYZseCysVni5f5n9aa/1WtViXaFYLBQTbSwr5
vEu60wYmzvyN7xhQlMM4EywshIyBwKmKFxIE5Jf0t6N9fE91Mo2/96Nuiz1Sz2Hh+2/TyGoP0ygh
m8+My6kssY7uwv0jN8lLjjp74tekJk5MDcA7YZJo4tO0csQtaDkaMLbrFYtiaP2ZKFySMsi6lZdn
XtuE10JsLQBThQrO+C3YpaEF4M5ew5uIFuUDdU4TquI2VKfEGpZxffqLzvjpPHHQ9IL9YXTunmVr
hek50Y9Cb447xZF/HlBowMGsqyeTMCeCpux6SKY5zRZSLRUdYQezoeavYWUYgUgRy4XrbaCDNUDN
NeHzKiHUlDHsMfIcD1/QNJ3+Kfepzk78oBtfNTHVuHwK6HXPqL0veXuxswYqukSpgCug+aIFTR7K
RnhfZOccHfH1h1KKvIIH6rwQbLYrIyo4mYQqsXXOvdo3/4OTCm9K0xAyDKM7bEpm5bJvHX0MB9ek
ZRoeOb+o84Rdkmixlt6QzAnkjswgioM1WPuo/r20u4RycCTFRODFJ2plNd/m7vNuDDQrWF45aX9k
o1JvvauyJVXGc9hIC9/8DMSvMJVufY0c9lDbQaT/TrSEGGq0RHxoH0h679v9BqpdoI9E+pXR4wKz
qNfezA2396y/Y3ocYiNBhhqfDoIqLqhJQYphoFks8d5G9GtR/jzA09pJblSfNB9yPAxji1PYfj+y
PNdMYrw1IrMeg+A2AL7eKGhsmXA+wi7qa/l+Xs7xYuYPyb3zpgs0I+Aw+mYw7L68Tld47qCMBlMC
nfELvMkaaGQ4zU5MUCQzOQ5RGY71KZwvYi4ifX44718KgvpUDic4iAaSRZTGwgZUu5RnMDxsuU54
gco8WkHNu5sjmKDZl/u+fKiHrlrQKN10n04yBt8Ts8H+bgZoxC3YDOu+FE8CH6oOX18oFXcRc7Se
5ROhW1NplD5Ak+mcrZgUXvmKW/Is7geZI6/B77UVqnG3F+Q3ADz40RXtGusUQIhE/okvR6aRN9Fv
GDrbcHkckXK2KhC8uH6qpuiOfarGJeqgNBcYCrhduf58li9MZlBsffzYF/nt3kPJoCZoUTNvnTy+
1OHceYqblkhli6cNTeU2VZ2MppIxcH66l190m/cJnLflMNmu5RpUX1LomP87d4IvtTUtjN7++oGQ
gDtA0P/TXhgAbUAV/MuYjE85pXz2eaJ1hWrNPjEsPdd8COGsOVuUS+xaG5nj00MH/mSSVxtuL6Dg
CXMsyOvA2ZZ8xxCotJ6dvYo25xPocabFUI2jo87V6bXc6+L1IqCHL2qz9q08kTuQp41kzJmk9SrV
VFUva4Ooo5jPpmd1x2pxuG24OTF3FtAsSTrEqavUM89dpxsbs58v5tUbzfIrFLALxrySaQLmD667
IzRhYNPM59+a01MbUiOappZAo7u9F3S23GSo82N78K0zHJAxUY/HGdZqThJ28+Fbb89sYcrAUldK
SGtce+V1CmE8XuG+UdBBOkLKKb5ENJHgiItDjaC67RFpW/1p9R1JcYIwiNt3vZ0ATQbJfjTPeEmi
Y5tqXwmJAuC1pfTJAW+bSCCcIgKrmfEtppnQ/FQXVE6tQ3cFek02zo+cbxcmHI7DrdP975JOVvWW
4M3jeGXLPLMnrM9/Khh53Qi7C2QgS7v/Pf6m/ewksAEv/Cf82w8qRUmXEReKFKGFEa93lrgkZTRF
k+pWOYodLEceIs5OZZADvzrMc+M852Vt1RIPq3oLlrECVXE2GWfVjYObAK0ByMbTeGJmNoahc2rE
T3/Z4ilIAz307K6FBC/eC6toKtU1Cd+tns2RaiBd+3dRySepivsVeyg14XWQAAS+jpcyht0stnmk
YWp+LToIBLwP53b8ck7SIw2EY2NRJxsFq5cT7ZuGhiJjvw9L2CaW7u/g9nJEIngc1uHxV1/CNn6J
iAzHsbc7nAVuSlPviQY5dUYssRRqhRJQa81d4nyAeDR8zSL8YqiSnhx0/QcfE+tHS6NlpYMtZhc0
PBi67jwwCWOKacmBi3b/QW3MYG5tZo7ifoDN/97OsGNEN2ccEgumxX6chNyMpRSlz9HyySkKqiZj
lhRJYIwPtYcrpwVCuOIcEf8t4XYIr8I3HAXuy2zUPNZyT44aBl6Db97LZomK8azZjUnHvh7lIjZe
po6abbh5t3wT8M+Itp3mZjk6kOkNNyd3KhU0BP1fRBIb4LocTNiKHP+kvXae2M+OBhXzvzCdiCvx
o7osSM9qqcFDGN+J5chE2HOqg23UWD/Yez8eY+muowwawURQAJx2/uRGySEBpFLqpGQnOc3IUCHX
g3LCJZTbx5O3aZB1y6CDOJ2Ko464mpEG8BMIO5z0SQO8mjzOmJgTjbhtex3EWWroz9LSwTL7uzn8
sRsI7nxSShBez5NVtXNFnbQs6i3H2MTutfKhX7wdHI5sswtdnZOUX80cJuAsQabAvBaN/U+yzyJn
akQCk1FwIYMGmW19DaS93p/ANOgylySyYG36yyZ5LP8VYHXi3uHrFE9pauxdssfX48OdfUnaeq3k
mLWC7gY9fUitr2t7mmA3UlJSn0uyWQwvUf8MIebktqbYPYG2/nS+yOCMFmz6ZKf7cAyeUG65HvdB
vnBI4PT2AaXbPT+UbGBcvNOlgfw1uu+Obi+icrIoYXbjT11f3mZPhTW/8bvgC8nFSrjeIrkg0kXN
QzUsNuNSYb0eJsZPSRvjlkwoMyDKEx77Xh/XNzXsyrVIKm37VIRxB1Bm487ViTcOb1VKF49yh2dP
m0EcOBd3CR/kV3Tl6s1nri9QYjleMHETl0T636viHZ151Ta5TVAVRcQbZlSgBsgc5elNHXgO6ZQq
1e2uqQDBh5Te70Kjxk49Ra+1iGT7QD+5/MS5qx8nbnZATkOnM5n/lK2pdnt5nnNutwp74rlyTbMj
G9tNMvZtk2EbjHl61Nf8yIkzhOzLUsnXqB8z+hIBrr8cFhwProxImNOBE/+V36BypcXYOO0ls4e9
VtJEwTMm6PSLzTeavYihq56xjSTd4J62rEBAQ0Rtx0Zi/7kvRiEI+FL9DaiUE7GO6Y89dphjzlcA
gYfWPDMJRSYiGdNI9e3jQRLxTUSi6YEb+12KKNflDRdbVJ4wrdYjy4eEvGCxS58M6TxdBBY71ghR
YQWSxwt18avDjvBiusKIfwYK5SId0zjiyz1nmIuq/usiRG9ZiivHBSHb4BQ3dMQlwDzVu0I4i+Rj
heGEixifJlgepCIER4rjr0RTkjnU0HFjDuuW/aNhRkNNLsgVq6P+e97je11YeLvSEgc5iERUrRN4
1JdR1J0vqeu1/MuOwC++sRIbSc52UUGn40BW+K9rhzjE0+Ck64E/HmxbSUhbzKpUzPDlIlXLgk5T
gZKQZnoPgmA3G0370FuY89xkUxurOikfQWqavAavDPWzJnXcUdd7LQOcUNztfeo0knd5pWozZb+p
a/UWhdyufmmmB+lPhU9Mqm1Ufq2oaprCJX/074VZy/8wawXELE2QevWmJaeE8vrOEE1L+QBtPxJW
wlvKIYsoQHqU5zkvwfVgtLTwAYnFDokyw0M3nIPYqNMxWFQvV2lqTdyP0XaGVOiyHH2l3S3zKLWw
7d2OFjIzQiGczfqPc3C1JqTrjQ1ulIapwYIXNwxhgLsiXCoZRzWYEqNZ66m8Dx/kz3cvWCQ1GQnP
ufVszCcyTCkv2+JA3uh9dBB1RyjUFeQHMoP5EvmP4IlSROZmC7gGuZPeUrM3mWtCYZ2frpkdnvGh
lLxp+QQ+j4PKdo5ww0yORcngSY9+omR1CudR516EuoF/dKNqrvSMWwZ1t2SJrkJ7g2TUfZFMyj9b
FrbAw/y6bk5WgVoNVwS/KwgnOUJqO6rvpb/1FmfN759TdndeHMt/UjqlavKIPU+F1tSin+T/iLNB
Q8PcV0sHOjByLkPHPwE0we1osJTmRJaSh762SdL8wdWIXCtPB5SHf+QBGBvI8hfot4A7BQGOvzwq
W66fLUx9aOHB0Tw4K/asIMKrJGqvIIT5Tv1HhQVb0XwW7X+v1cteiNbIORp4g/C9XHExEZd55Acm
MacO51seWc5nIHr3nkoqRBSIetjk/tkMS9v2RV84CBMgMmTuowxdwy+VZ+U2Oq/mD27OZ5LCuDz9
yTv0J4Ker8b+bMKyHZbpreYj89BJf+udyX3iCljEVlROYUR5QgmysEy6bT/+xFueue7M/wboCvg0
Z8h2bZuHja5l7vEukkPYhlcySUp4qSKWoQP5DCdGgQjwoUkOByWmT125tzglGd4n/aT581teeNki
2WVRrJRXG3BmvyLP27wYfwRaZuNua6GYyjofTQggyvf4wR9gmqzcfGYDXfniW3H7UHyNbOCr3bCK
Ca1favOQboUTZoo8T20EDYfukQ+rbU5vBgFBI/enTiqGpmG1mxC70ll+F0b37sAcuOcJsJjRQaEK
JdeBHfCIrCcPQd1V3sTtDUY44E8T33zcQuT2mKMfdYpJchbRrIzhzNbVxDo5NtUbBgXnyrBWO+Ez
gWeuXqzSRTx4ejBZ9aS8hmAj+1T7Y+ziJc+lxnOnvoeMO+lyeJZucq0QTreRBn2hhlUyHrcTgTq3
17tOnjdSCECfumWQdkXQGHDgo7QiyOLgWD3s0wxML65Vmqdp3rAdx82+OI9p4aze1YStbHhDRiYv
pj9TMGIIxhEzyWH+jD4/EOiXdlntQsYqNwHKy8HYgTUlSmSdPilOmzUofcvibpWFPpGyDorL+9DX
6yP0n88A8FABfpk3EpCEB40ypkWBXslQRikdVX4inCIXmzKKu/Va+XZJXcl5oabaWOViIwVm+3kR
ELSL6JwhOSHKU0UKZjgvritlFpAkcY3tvH5KEkLu5miAS8Z25y9gAcEhl0terbYgjt5bkg3HHsHa
jkMeluIQ+l+FFeszdNoIByF2JK+og8ViRn2IjdeDv4397i4D5BpoxxMewlZ7AJ90ZEB876j4YRJ4
bL0NSe7yox0JBUnkjQQxOXYvKQPVlEC34ONZwrlkuBAWBUFsI3V191tv1Biz7fN81lGYBwp2DM3i
rmV4OwULlxszs4IymtLPVo69FEzm2f4AQ+3kJx18HKIL1uQ7GCGqorSpsG166nX+wWvLfNCNIlMJ
boObWA5sUEnRzU/6Q19bd4odp0+cu1WpE1gEKoVmlbBLMDwObfFurqcReLCb2N57wISE2FcTEQIl
UDqUbbpUv87FpJBwPblB4cmo/NcpeBA0YYUoiAHARnkVPo1UvZv9YLHRHM8VlH/2fxgAOAcefG4a
W7/e6AzKNfzs3n+vkXAYxLWejSRhav4iEXVuodD6SR/43FhEWkXYT+d5JMWaL4kaAMCOjf3Zgbkx
tTBYYjKjr2NrZGRlcqkq8YM7uIU7datqo5thJCNMyHGED8GEigNTOC6ApjZyukm6jWVOXDQnVVxq
jL5Kk8F6TqLJjS3sWvdf7uCcmWuZF1I1Wv+mGoH8/UAxfQqJORofZ/Xm19nIYMVsY3bETXFTcd0o
qhxK3qTMn1MXJgo2olzFezL/h8FL4IC0jA1ECe83UaYvuUcfyvGsFblekCLS0BhZV1o2VE/tIe8+
HQ1HY+wiGb2eCh64Jw2B0CEbSAmGyPZmMTjCYHOnrFRI1PoErD2Bfm4vYpumZ2YvsA6PB+xwOjrb
KrJShIt/pdLzviq3iRdCCnO4LJf+F7v4FU44c9GnmFqUxnXgKvyy3Jr46sggWbAVCyr6MHhktib7
R1sitJyqirFw368LoMuVFDhomIy7YrJomLZWj8FOkXvtUshoyMZ8rMSnyanlR8HqVc3vY+XJw+Cx
MywEhZtF1+4FBV52Etp1/VloTw3TE/nV3UKwJPZUPGQd1h+VxFiHiyAZN6mB5USulKus/ooqjBU/
Opq6K5c4lunYw1LbSSNASEJuncONRrfinqd8Rhko39wT9KgD/oUiNaSb+SNKbwxDH0yiI/8FS/WY
Tpd6rAF1MuHjyUZDOtIaLDzUB1FN0muEL5m70GFP+3vHoPnPqk3q719szcp0ooaUM2Wh/l5dDKqp
rMoN3waOboiGjwwGwBDv1YMwf8/G0NRsFRhM+tIS8RO6rMUqiLz0WaL1Esm8TVsff52Q9F3P2BKw
/VeGvDOXB2zmJkPj7iLeVv+5jKEjEn9QE6JYobdOHVIJbnjTTZitPg/Njw2HUGSxrqMqEbGDWJ63
BHYOkMD2jFfjrDcnM1Ru16k5GdqAxg3oGhgzOmvlByyzogdnPmjt1i9IuvUt1Fednsz8UJx3XXqE
wceouCwqeUUR4Xa65CUzmB1zho7DOZGVurlfhRTGrRccwwZiPyZMn2etSaGCHOyxphcKOHyZmH8S
G7RYUSDsvnx0ZSx1JitEqi4fMMY1ECqtvej0oWrdz+A03jnHAp7iqlOkBT6l7d49EXef9dvKYZAq
F0cSRBo2acT2fmedUXMyIlab4UTy5RDM/9VCJnHofhELMK37Xo6OgSvgOorwo2oXTRO4/zlgOAxC
N1BHxn5o7VyrcnBez/tSmvmOaU396nwiWstVZ0CFvJ5XHWIMSGl59Ab5KlbHB6NHYG7L1H3RxirC
4nhYINEX5dC8IF+ndEJAtC6Y83gnQomblefbwdq0qkhnM2undiSCbT4i1Zx1gaNzeZQzCyfaMPu9
IcZwmRts0+/gy0fqKuv2aOlzQtD5MN2e8bpEYPTK0/QFvjohFNID9Gbqnr7/XM9YTFCPzEjMDwpw
Vg72o5ljGbSIcDZS0ldtnHGqV3Ipi0JFki6kp1pFCaZYvhNMKpeP1AcezaO2B/Z0BXo+WLO6tz6K
6I8aZsGYBPNSDIb13XVg6P63hGt2+nPujUIsM+fzl5PePxy52H8X2Pp/vsd52rExXPN/nls1yhww
sR+SNyOvC0CSLIiXyCccL9aPuGD7VF11WjmBeLwhbE8qWrFrKmyOx+QKsPfZqv9/cxn9RuiP3W7W
IO0ydE8pq+t7BRf9YywwtdpSgMxpP3mcL1HzQ/YyNMr5x9W0Q0YkbXbS68ZXio5EBar6LmyZ2EV6
ghTUDk/6iSvNKU2MsBs+qIUo4MjRtPri3Nq4knX2e5Gt3Hvt2zj2B/n7jCFYaUTEEnWAUxKHjuo5
ulalsHkuveO1BnjAxZ8YGTfDQeQ3QRbYxPFC3DVJCEvZ6+qxAYUPVnZ0/KOVjR7x3hjY6n4vu322
M/Ofg8RWK6D9ersjnIdz1MIBUFCuFy5Xs+QKoU8e+uQ2WM+199GP1qfi0cyJU+Klia+qBxs8+wkR
g0eXh9aIJUlDNSax288fDbikHn0zcDX9e/ODNPL4/Ay3VRGMXkJMMBiyeM5xJQQxursWQi1f0M95
Mtr3YfRY5L+WwRD2pRggI+P7xykLSavbxDVnOhXMn54cTF+EoVteOZ9f8ZNTmWal0BgXmGs4Yxth
kqbldvu1+oZsYnPZfqmMiMheSHJcVrBjP5GaLEbFW0+1qn2oDsSUF+yuJoROU0hZhFMHddnoLWJ5
xpDzp2ocGP5ynDe0LHP2kNn+DAD2ckvigB7NvtKh362VyEQYCCrZG5W5ift5BOcflSQ72xC/qsUL
4ibOSciiwpZSFLpEyQhgBo0sQIC2gORnxdAMSnu/uADpmejpg2bSz0ofXEjw3keCYrehj6G4fbzZ
jawhngFqwzvaRO3cUjNUkMnB73v/W1CgBOGUb+xJ5YhFsoYnFIQloPfBLVg9HTZmEGRDmA0fqagp
HJ9/KqqnDONx8GLNmNzWpxFzh+imtX0iKsPMxZAVx5Si8nK8Y16nvmMZgWgNW8bD2FNv3EWy/y4l
iHUPBqTbsRGIvi3i5HKp7Hd+NlLaF94Hh0jgVM0VNgc0LK+fyZ1wr81UoMU0FchanVgCI1puyXr2
eHO5utNPaJMFWoEtcLeQh6AJLbLPi4mhX/0aWrEF/3BiQQJTN4hGuxAU14si3S4X3f/GfMW68TzC
zfI/eP9g8exD9/3t9r2sw7/irJT562BFxpJvdLUcpQckT6I6Y8HAKRHAiB3tPIFIZcDFO8O8cJ7r
NtTXHPTkqW6n77OGL3z4tc94/VWYSHYrnWzNOLz5G57I2n4GIH+7k2Y6F9GwTND772MTGcyJGRyy
nVYYTjTfwQPm9v0uRINXOfWhwGBr8CT/bW6zkjNTBM9csy3jQVcxvbZJ82Bgn8vSNozNrEjpJ76w
Lhns9VqsaBADA1Ho5QQHnpRocb3DMZcqkvP4pU3HhNo+hcbfDQ2mNgKu6/qiChNY9K2CoFFBwJYP
ZNOU1/vBGPdRJ58wVogr1G2M3ZhmW7+jjxSNYWUlL7Iv40EHtbsnn8k2HoDhtOSTkWSPQmpxUR/S
cCVGdY+cUaneegYFQWXPjirmE84D9tOTm3wqiP9v7928FUSCJTiA1wMwVaesLqFFpQIiA93+cQKe
NqtSyDZ6lD5B/bFQLX97YQ/3Z83bq496WDTh5YAHkL5m2VcV7lEB3stQ9361QcczxlQydW9211th
iVqa11J6APvgnz6pMefLHMW/zZlgxy+xtbUEEhhwI+GZw1FLybwL8yu2qKanPCzVjbWHtyINqDeu
9Lxzsha1vUqr5LGp6Od9SHDUFgPw6LasftVpuC/b+PCuWkiTsB4SR7krg0NKUWGThLjhQyhGWMV1
ohiNhKuZNcqZcdWwI0LwiwGczt+av/VF3WhyF8RUUxUX8nPnLVLxmnfNkdEDA3XOVuzQ1rfkn+wg
RxN4+GLCXk+v91HRh6zTvPmZdIth+kzWuGYrSjkbYbrlEr5i4cogZ0D+qM6HRJvEWYNncawqqtfL
MHnwZLvGBkZ+B2isqEArpajX81W6ZwzI5P5RfGuNM1Qp8+nlhHhgGFwkQJ299ZZ39aApfutEUoJ3
jsG5GD4XC3V4Zx2AldX7eXypyBZokPHrhDcjjy5KOb/hPmemX+w28K5xHfP7h6nRSbVaP8Po+6a+
OYp4TlFYv+KpYZ8IVUQhK6BuHiSY0xpepz37QLjD8yiB2eMhGGMzMAdXke85Yh6vKIDJqukTJ6Nb
2gURpp6GnJIjt1b+q5bS8BQ+cvU2mAaRBriPVcr/zSs8F9jUpJ+hGscpdK0u8mz1GOgZ9/K3Yr9w
i6E92LoGiPcALm4J9Rgc5s0kIKAlYqm08CEO7mOsYHSJcfc4M01FQ5S02euWTC440BEgM7iFNxny
yD5HwYy8IlKfs2aY4d5TLG2Y66O/QilEStXyu6P+AgT/ycJ+27hXwiBOfC2hR57fF8ZSCfI9kCRI
1GeUK3poynMxaFLxTPTtz+n1OC4v3BfxUebISQ4xkBTlBIEleqRYjibBrr2h9REYV5vC1ugWvxn+
LFevyi9FHVzhv/Rw6OF/VDalW2B8SoDRdprhniuCdiFrTr2fdpMTUH22xNDexVTR4wLZ5vKmHZYi
3il5cH4UZUUyoQwqvrgUXEMqyuSUVJeUDoTPPWMHWaVFLfp6yTHbe/+zOyl+GK8R2AScWikEYwoJ
fz84pY8/ESA5t7dsKPLWE4e3pJeDDy40q8OB1eRhZ39G0abuDaXbZsZGhiU4BovgBzaNvO710mvo
Yd4AjqYzPL+Hob7MegoLRpeQDb72RS3J0gHtTx9trf1zwwvukvwnH/nFswxYLTNKufAPKWR7QQfo
90n9JmpP0FZLSSlWyLMmVLbQYx8zRuVXcgL3C29t3OuYbS8/bv7VBEglVvyRskqiFSHFmBgCO2uL
HZRB2+Ovsyc4vwYgsasD+ZKBZTRbRmSNLAcCB60igYIMwVSISabJpYxhPK6S9nbkFQL7wsPWR63B
6P8odOvNFPYcc/L/KQ0JhZP0n5t0TvUVMYo+QaEwHT+gELoT/27Il11w/HaKbhccSn8KyWdBm4FO
LQ75ybtXG+KLRGC6uWqyhXvx0hppoLnQpH/CnWh7lyWGiT4ko/9n6GHLmVRQAnApJKkofHP/chSE
tntSQ7a5at2QBoEBuuUnEN9dUP3eAIKDpsf9ZlSe7Nof1fumKu2qaufTjGbDrIjhggZ3Qs+ix99M
p2/Fa6peABltKSMSmmVRLm13J3r/C7VGMLTwkT3eFx2U/4FZWg4RAhw6lGMDQu6OU+0NVl0Eace/
yv3f+obGScPVB9McSjSqpchS/D7rzfGaEwzwLoIOktA8mPGvgfSL5ca9Ep48hs0pOQs4Ne+j74V6
aZX/mAqdvZ8nf9P/15YUfRfn+OkRgD8z/ky9D+p/cacjbnvYqKgixLIEQvM15kZqdyNk+M2D1+mI
t5Y5WcLzc/X2mxMLGIY7WcynQRMT8m89AIrSBXPlV6w1CU76Oq6ykBQlM2rnfsyAM4vbs15UubNi
v8lX2Dl8FnW77Lcr/nK5wpAzpgk8NHHE08PEzfyZNEGeQI3H6tlf4wLWFmHcLUXaKRWe+rQDElge
r215RYII23jdYdv24PiRGMfrMoM/cCwPvgm/YiYTDvzCjr1fS4uz+vUNTciwElC9xjqqsHr23VQA
CXSsakNm7ecVjl0cfk++K/jwEoZPebVY7HOkevzBoESuB1WBJq4gsQQbok1RBJSOewOBkyJ325dV
WlLQjf0bbHpMUhbMUd5i+gQPlhDpdk3p63vLKkIY872Kceg4H7DIjD+J+TexU0efK/BCOdiLlwzj
vhs6lJbCcdwFxheOLPi36Cd3mOahZ/CO83mwCRu2u95DdjquG5Ju9NMvAp4ZBVjB2GsU1YV5DPV/
Zj6PqS18txjOlmcOL3TiGDMUrVugOJUzAl5txMLBhdtqqvqBl+aRnt04uCQ+lC1LRR6kGb+RE700
W1449r0MQNh6xcuDq2rHj4ZFOAeSHLP3CILcgAVRh+Jh4DpGKoAmmAyVZ/a1dMVbu5HU5tPaksga
gBLyo/b/HDLeGEk0utBpoDF3QtrXGTNVqe/Z416Gdj9d+DqTuIcsMExnSKfCRYqiaa6IijMm8Opm
9aq1vdnz7JDgtEB6si0oKSJ/dRQi4S/0AZVD1W1HeRBO4LMJ+oHFosAWWtH1MDP7BxNvIPFRe72N
vLUwZG4ovPhx+qLMrfXLL7v/tPvAM68iAwKa0AEMKX2Wkm77dgJT4mjDw2ySBaxbRG/QUg/7lscW
Xr3Dkv/Na4tqyN4BqKecRiIowJ0QjZ5MHl4bxuUwTiWjcFonX9eSDMb1WY5EIIE+JriyOotq3nIS
ho2h8Wf0Oal9nDTxVwFbklFxX/v/bwQKhFcdTnfp3qc43q6ZwuuleOBhQpOoKKB8790uzWOyELbi
MMnpt4SVcgVVM0x+Hlx6uroECDlsptsuEnsbWeXVTWUG6tedlSb31UY1ZBn6UxFy0WGkHw3yLwBu
4JPuAYmVmntMBdA2v02DpDBtO8l19bqH4rlcU7sTlZRsfCWQCy5UhvX6AVWhFVjais/bEnqh83Ck
BZC3cwPMoaw4XGNtAkg+B1v4s0M7ukJKsHcIr1uabqrhD7rQ30BvSUPUVaHmyzdAZp1q4Tisg5VK
KWbKkYn6g5HaiIVepityW/qQKKomcUHsdoUbaJczT9gHrLXJpGjwtv0gUygKHpDNV3VHqKjlCeXh
sqLRvPoAESn3wvFDLlhY0O7NdesuZ7ZS1B9DWAtXy0vo5swn0m9SmNwvkkV8F9IpSdtkGh2mra1e
xpOLSIBFjoTmenXqWuO4ex9ODI54PclXr6E6csQrCj0o2dwQ3KOAJPDQRAX+UmEvI6Qop3xpAM0F
xXzQLhDLfgYk+H6S5+byimZrZfXDSA6V1mlRp01BQmo4C/RBA87r1FrFtIJip+wSC7BHDk38oCLw
I/HUCUMSJrBo7iax/AK7r+QGhZzGgReKhyr9mjXr1sPbUwz+NgcBRfX1jfIHBcZHnSwNuakCbPbz
zzYYCzFpX83rTS1s4cQB0sD/4wssU/S92G2Jj/+dNRcjr9qAcDwrvnRy0bywBgAzaJFvsQmAmBKo
4jS7Zz9Xgfe3UMHMl4AtNjRDjFmGvzqRLOxyYDv/4wXZtJRsRy7hH4XbJ6qkxCVn7yL/TfLweQel
CGiO4FrkdsdTYWqSr02tw+hzRDWgUfUGeUiP4nGBmU8nBvHiyZ6DhU1hnmG7yuAMT7h4/xAlL1Um
4TBWDhmVHq4J7+c60VxsoD4qy0/d/Qz5+so1LGaBWf3OV9Dyq9yi2AQMn8pw37w2WOSJmRpXZllm
ecDaFE71MAXLp/LslZM37kx0e5TVhyS9eLUSAVrw/5UeX5FpX+mFp959+tSI30sCQBCpUE0cJdg9
yuuciHWjQum+KPDJB6kWKpEqoB2cmyUqV1wm3vG/UcErwJw0SNGxKD3nXQjY0s0YRJxt19DON3yn
BVi8L4IQeD/1aMGB6xGAl4GSibbeT74kiDta6Ibp9F1wJ3v11zmh/4GPvJjzkXuP0vuB13KAunrf
6Glgdjla9VdI59jOIixEKndCjV8Q31ysnJmJA81vxX6J17vtgEshvazTaNtBbzYH0TB3P6bfMB1h
RQY4tC5lv5OG1ELt2BDaYey+RTfvWLfsaq+Gg2UVrrmWt5YTO2RsKXGVUwyg7xDjrsL+EE+VeXBV
wGSOj7Noy7/dte/kqJw+F3e848ClH31i2yrxo3gbOuVzXdSB19HI/RicGNK7WkKPQcIlk7DZ2VVe
BdyZpKP5ulNPj6W1WEdWro4EmheGMKtBATBhtpVJXD3S/i+VFgRZJQ81Fez+vtyh8rtv7XKkqyoz
JXFUSGv1AsQ9zaXeCsq5doBVYoKSxJQIJroC0pZ7Zwrfm2XW+G3eOVG1J5aopSipH7zi6rU156ai
tftNP1PC4Cbjst6TyNZoXqx8gn3y4sn/OfcoLtyWNBwpqJZG4OM9Tjsv9gvXq/nGNsp1AXvoPiso
82ZtJdiIk3ryKFHOlecMFrUYs2rlRQ2p1oAIzSdn4t/iXdp36Ss5tI2MeCsVXQNM+r5VfnW5abjc
91ud0drsZauq6f2+Xx7ED7vvkLRS9mAABgJW17tN73JwRC7SRyiFspaafzgL+jRss4IU10HiLcWc
yhnMaUByGI8H9iit81XWRBfwn1v35CEnhzRUrKMmo5HrJpzz2sjxSJFA3iw8Dh0rMKM/BoRqdBJV
9ZqIx19vIKjX/Bc/VdgPuCCI19KyNs1/vfqHQjDvyAGGXz26xiIIaSKUotaWTGx7V+ug2kJn0uFj
DAVlsVGC3ToBGl3ZOhH8LW0rCfVJxSkKUH1MZW/Fmx39fqR+gsB+AsE7ZSnS+FhHpbxNNRMNukVQ
eGD7H/UO1sdZpguldnmPvjSGoZjQrx+4Pkr0pHZt/EsDDlUjb0XHzpLHOxnyjYAUhCjA+fFKlPtr
7RaLmZsMCjyrsBwnLTpWZWIUwAfOWXjNUjzGDvg1lftJdrrvGUIa85Z8DwJqWic5QlBY/svYwv3e
1DCKPoG8J++a5/7ZZKu2SYWNj1Kr6i2qFKB9AhH8Peg3JN9M2uYOV92jo99P9I+AXU02XygAwTaA
ydoJRQy3Q9yQTTaIaj5Y8q0UO7LULnmcOessdChxNlpEXRtiS/4XZpRdKDRKN4e9GR/CovcWiYhM
KZqQYiajeOxZDi/6++sXkjsYA9teCNPjpiP98JcAaEOjj3lwUlvjZXVz7zQj5k8/WV0xCTjKY7OK
wwM5Q7dify3A1zBFL7lqmjT/QKGSeeFYX7r+Q2/cxYPVIjrLVFYWdAvkDmhm8Z1jU8SPLRXfIdz0
M66X481tQ2zICRcc7/+dlgdPw3jeGK0jlEzjZ2qIZFcefLKvKH0H6tpi0lhft49bp0CZmh0zZa4q
EFGkjW4nIs69MPpMnNFBYAzDfyxpbfqhxXRtVptLFHmylJeCrhiaKbzV6ymwmZm8d+mUlMwoDc5H
5pfvjhA4fJVk/GwmuPkqxHNnuJzmcvU1PFRg8kKzq6gCWFQLHj0DoGFsKbbM6gmETjPWcKlbr2w1
kNShmi+7QOCKKY2Dj1/tG+1JA32ALf62djEV+SElwSHhoqah6Egz4fV6Uys5OfhKV9fXWwNkRXHg
EgT3pGzZJUUv3NO3yOs4obh3cBUv8CAZ8Ok3Aob4EACIcou5ld7R6Cww0oFuDv+ZMEaTM/0ds1sy
wwzPJohuZ1WEwgf8gMIU4N4pFke4nl79X7C0bEmoZTj4+ua3I8FgVZTVBz1jNeyBRTlfiI4q0VUH
lSZfWlMQFRViLq0SrDkNCggN/yMlkC73Lms9/3zNWv6U8HneavS0hNKlYbR0LoQVRh6xJ8AuJ0dI
a5h/rvrWr40DSuL0Y8TGjmVacSNSHWI4qB0o8tj5tFjP//ChJkf2+zljS9Yv5tBQrTRl48pkGcHe
4tnWucxLKbkjUg7d1LvpbnHYpWyGcpjqHDPQbonNkHEGzuuaNZQ8jM7HOJ7Q4wAD99RafW/ZboS5
pCUMP2V0iZiQU70IEHWOO3MaE/rfta4d1+ccv4oJN0TLPWFmCYziMB67ABBfnU5+kURM79sA6e7W
E9xEWMMKhmZ/VlwPdEIDX0e4/6anPQZ6BipgEk8pl72HAPosPOoS+FU1Y9MasP+Drqyl8bH0qOro
y+JL0QuuVHvkoN7hTVOWsP2f9VvPdafzuwqTjyFtRj4X316bW07Yibe8axEUMoNf3gaOsEeGjrMh
0/obxuCNNOboKE7OrehxIOxhES1vNM3n1snzOkOp/n2gSOWU7PTXZIA9rk0jRBOYqVSGalGaz490
0XMBZ5gYut+ied9b6IxDf6dET6uw/gV8+wuY3oBzhvpwpI7gUpP+ZHUHtK/ATkxnQwbSbBy0oyeC
R1sYlPZfjD73kx1i2ByhLO7zuKCpLGwOofZuJ3CF/lb3/MJi5dFS00cHX9m7iqFNKWI2Q2u49acn
zsn74zHMZChlwq3h+SAbtmSVGC8ZJamKt0udYQZbuvw7oHwdf68Ftg+jaObilMfvXK/FOpcd78u/
osJIEOANFfyJnjGAV4VFNruGDulKaFjRfRa+5iATkRuVQOnQFR1E4i8nyUp6tF0T/cGcaDyCGqFT
2Ha7Bu2Jnixp5f9cEmitI3/h5kUKa5UuPOZvBlj0W1hmZ4ZuTgZehPfmzyuiQfvxZx1uI37c7uAh
vj5rHYKP/pkgk60OEaoG2QBkXUZ3RNfm1QgGluAYaaw1AYtRKSa4+nM2PoPIfr9+akiCXlhX7oc9
TVK31l5Ro0vXJuRfFd6iKbiTeVRWEY4rDVWzpKTSBuW5orffB4vaO9a7A2nFpva+nBDSdD9yw5jX
W5aLgSm3zLc5jPKVH/ZLryVr74AtVs1ajUBFn4M/4BF1sJRwQk4DIXBvnbhpTmShwCiQoPx6zmRR
zOiuNmZ+fgrnJhmt0ddG3ODGvga8o2g2V4iJhVjg28zp5E4CXow7AoF+sSqZfbbBH5tQIvMwCYDB
8DFE6WQofMQ41svlw7FQXrfrWa1iqqBtLpBjtOdihbtskY2QmGTjilqVJvoZj209DipC0uf/IB59
PGNHi7gGmEldkSxtjcRCYhYPdtMX5pzkldjbuJGKSGhvgpcWfhXisvBuPeyhqrD0E/ICX/+ZyAub
4Kpa69Zf0rW/x+exqMAWA80C7a66/Ttb5X2dfWGjQRHwj84O2dqNVmouLUh4lujASfbjAoyJOiIv
fDCTd3LyzcVCwpRF/o7ozP3Zthqnezh2PAEKB7QOoirZpmZo9E1jLzMlJKe6cmP3LuU2BsJkER/q
V5Efq2fV/mvs6iSN5BC+c0c/eM3Nq8IepuW368XX/App/h6+oCZSGN3BVUYNg4TimMMNr5KZtKFd
fJ1DLmFGMpyMn9c+5Nxt9+3sOim+Hwy+isG6BR+6hFo9MN9HU7AgN3WnKgllpzRou4PEPRmOFZE2
3ukzb7FLSyKKt7B8wQOC2sUWKsuAabX2eiEBB1dvXe9f0aSimhDEUEi5KSaWz5dpSiV7KizFU/0h
FNs/Bo0MQDZlvmktmbLndo4l0GgawGUlZhOTNMxGcs6ASdlH945OOhfZOiF9Kzrbr9oBA4MjN+9w
qkYyeCIths1+191CJEDqjPVVaPzzta/4ghiTIoo3xKPtlNxo9Uaf8aqPlzNwVi7wJhkfAgvXYCkP
5Tpc7UGNvKBDzurJ/0fys2RZGKr6kAtJ8ePxdGoSMmDwffMdn9dCzjVAJKGVGMRAEWrYT/EFwVSv
cdgbfIdLolZYxsGRkcyHzF4bSP5Dz8VjXzUipVO0GBKQiXSRed+fbI5qagb+uDLTSKJ/2AfewT3a
kcWTyNDdzRIoWMReD5nAzLYjLQXO+qNA/REkG+WGntKOpiAIZOq++ZnNn/HLXZjrPiXZIB4drzLb
uduzY3WPTztfd/ParBkkqgB5jiebA2gzeUuqHhr32rLbeZV3rEeZMUryYhP2GqCZkOidw71AdSMR
o4kzedubs4SR9U5fX/lC2mnzhwyRKFg3+3AsyeytJYg9eEfoXvwVJNn1jIAiIC7jOXfCIPYUdbnH
fO3W/FmlsesapRsjY4xYn5hLEZnHfFpqzsXONrhJIh265roImOJKN8hd3Uc+PGfdFED7WN/79fcu
8CXfn1mA00WQvnGpsWk/ArQFu7Xr87bOsWF5c4s9byCUrA2HSew+Lwwmcsndg40W944yKdqRKH8l
QnYA69XnPfd3LXlkV50Vji6Y8KzoPakA6GRB/nEUXL+UcpR+AR9lNZbgecVLIH6FSjLLMyTyXL2v
y+8AeTEOkSekYJxJz2AcjlmiNEp5NPjg4yoAul/OZO9W2oNAl6Yojyy4yP1rA1xfX4q2XLBwUHp/
gzAu38XSClMTu24JWnhvomtqzIRpF+t4J/LdQ3jJehNJw2OQKOeRHUx16dgSHhBrLtobo7pW2rSI
8rJRJ8hTJiH61MI6g3V05I33yI/VGRHgADMFxJMwGFe+b8Zqqzgfrq4aegdAOpa/sVovHnNhr+y0
CMMyCYt1GjA2fQQsxZwDSkvwHXnGDbzwrfSV6AqK4sNlJbYlwYoqrIIx3Kl0INLBuT/fID21T2hw
iDhGd7sjZDh6616AWTVwqOAN9SZTVE2Krg784PCaAavMm/MNYBTQFGhQwR55/kue7djZgrS05qJA
h/FrLcCZ1aGl21z3wNPTorytkcTpMcR9wC9+k36kmQ/uLFJnia02++UmheKEvLHFdOXJ5BDeheuJ
yE7gsUQvbk4lWZNlnYED0jv6n9hJhmyLl+6C0HkIK9oNT1FFZzz63jF8fMZMIYw1bcykAHLtVtNG
qZ6lGaCD8xxXl5CbdnhczkFnNHiWCHaEUTs9kVdAB4TatmdW6GidF39dkTn83VLpLAW6tTh5dJ+d
WXkjutEkzy1QLbX+8APtV6u47ClJwmeZ/tqoJVU4foJUQMqQ998N1ZXHP8KoHCjEAvUsfuBU3z5R
Okf8wLYvKHANjZccs/AmmMb8J2XrIiysusRxm/a0TrfcSy7bB/D/65G2Uw4qoAMVVa62ieoSEEg0
cqbF5kswyMLggOtTBFCtfqFplJcSK040Ibt0gkq4W+1DLr9M19ZeQL5HLvqWyiK5Oa6slRWJbNPW
dlEEVsY3eo7rxR9KYSbGc7rjDf2vbXhJ9UKmP5hV4F4MgjqzrRA4nSe5fz9ZQ0YXDmmO27Ym9ner
q9viOYxUtG/roEnR3OtozopT4nD0idH2Unil7M+9301cyLbILURCA5CXLxLStqRsYfV9Q60woex2
BUIeHsoiqt2rMisH1GyT3gHQQvoLK7mvLWWF3ZSyabuNycwooNTrdsbXTav6XJ/e0cADQvNxJ+8B
hZ9CT26f/PsfGKvgd90UMV96Tmg69jgz4GvuEiSjvqS0UYM5efWXBDmRY/r79M7tWgknBryHyTnV
2je6jgmHgubqepjMjg0zen2bkO4QqvS2w9NfUjR/Lso/SDdXxogNyVdri08FjqZuE2krIYp/5zHw
BcsqrdcHb2Is273x20/U6qRW3hRdTcp7azghG5zjIc1MAvivbtnM6htqSA9nCYVa6nj0RN1bz30J
h/2Dkfwidnk6pWVH0b9yo7K8icoZeIKpctBLOOcY5WyDOTvbWjbZj/g2Z9qTs1geXh0vhBkLQDK1
x3W1ZsSLZBlzVMNESCo39+LYloq86wIp4QN1YyOmf3M+KFel4/q2LG/gmztaPprN0mHC7CPXz3R4
7gWotfBq7pkAWsdCuCiLfJ6e8JrGMbanVmTZXDVwBGvhqowGeaf1cTriEiwCi1YEBz7HHuHW1tAi
kCuDQuxlaJLZMWPMWF+3Z1apBzTTu01cdTDZw3DI5wFPoJ5ix+rhQpW/J69VlOSr/jUZZeUpEiq9
4WFhcJNQ2is9snb2R2nwJWsSvsoah6RGCIWMZkynKVEfVNjMuUsOIUcRwUbyWz6/3wnqNi1Wax+3
Tenz96AMS+sXETFU9Z/uDSfzj07Ysxt9zoN28O2A1IARJirbIymKkfi+0EcY0vnSoa1BJCHlV2hH
NnwJMfOPddIjg618ElnpNzQLJSwGMbLJsaJojLN9gYcp0Y0KfJ/3epcQrBBBiWpNQMLFJuySPHzv
TmuUhX+OV6lPlAPYVLXxHbKunHZIpAV1N2hpd2jEOHk715dJFK31Kk5+TY37d5bTvck2YUS/jXpl
bo3KZdmKDYSDVOFym1QV3sayTqhywBq77T5n1mH8Bd7cI/Wgt4ghqRkkakCF3rmeAclwjQIk1IXV
a0OEL44iz8zWv4npXdfRcGqfANqS2iqAXIm+stxFbtdUh9h0FTo6zXxYaJLPUunWtZWZfEmIruuM
RK6azBt7BghIc5KNN+sK5PRWddGTcQiEszNsyHWcecCf5qZ3eMmDnlbGSRcQaJAJTUWD9l2rifMK
+16xvRI6Ay645gCcUP56ZJ01mM01IfowfqHMq0q3EIwUX5753/sJFQCz0/Q18v6LKWSpFruNJC3+
4uOBUI/eNeiU+meiflRLs+eNi6C9TK9ArNS7pW7FNsgFSbnBmfFfE7p6bC8qYfO3qHiSpO5qAcOv
27rKv4Sn9MhYHHqWxKNVSFUSFQclGcUMu4K2osh6LppWtOcQrUIMgVLFqvDHmCsFhtZ6IOc6Rux1
wROaryJRfW3FIdkMjYhYjzlM4kWpFEYfhr5+UtUGOGiFa5ak8/q70LsEpmfrrzauLXGmXUNTQNd5
yx+P7nBaDiGmdiosMF6Cy/5wPDWd9WScdZ/WeHrNc14ikrccQ8+pg0Cx+nZ4W3qbdn+gg2bcsNMm
+1pacvxH4dazXBTHKUmD9s+H5n9HWQbuqWCZLCnJA5FcrbCtUStMMh93BEAaXBbA1Pz/oeKXNTQZ
cTC31LQaMTuPXedDlFU0NOLEuEOb09nQeVc735ejd5GzV4gu3WDXqMiiDzuwf5NI8RPp5OWK+td5
eo20qmlbJ28UK4gd9cbwcCkaqxhTD+bRhdvliFXDQVaZWDfiFkvhOSNlV6Wbs/F1l2t/L7DT8Ty/
Yds+gUn49Yd3hG9BrX9NfP18OkXWtW82FgbUc5zrtlQc4WJP3Y//DkAIRAKuTAy3Ofb5j8sE2mzf
szXcy8lKYThadtTEdV+xGlNrvKQRrsyMCv05fR/xZ1S1Vy8H8cVvbb5ZTQeQ57Hd3EZt0kmF5JfU
hyINHUMOIKki6bqV8Zli1154J8yrj+kYtioa9FWBZQYQDyoF1+iIM8phkT9etSyDDo9XgJEJ7TOC
qd+XLQCKreP7D8cOIfVgfi0TtRzM3vZGI55nV3BK6DKl+88diy8bL0PH1pgLJcx0tZRbxsTvvWQR
qTyOZYlWk40KfsLQUAM99eu1B/nVwsp6B2ZuNhQhvgCH50XbJ3dQra8sEftAfD3xxGaXYQYFBW4m
r8+1ynCieZNHlzePQTXgyZT7c82+HQAqLSBAr1bhtIdYpG+YIk8gHS63jrRkSsbvnb/20yWH59HV
52X/znPkaBHwTtmi45WaiSXwPsqWeWxQsmA9xMOEjEuIFTQLoVMjNskBgXcAloqva7M6nAo2a1Lq
lxo5svf1Iaxj71EA+JXqfAejfs/piscCOaJ5RcTm2L5CucyNJTyeDWr19q37sEzvuTkes/OyjiAa
+DRpYd6bGfVrltRc7Wr1fOETdaU5dXPiZRm9cArTLhZpJ8+CbzYo713B2+vSTp/cSGHUbOA+nYcF
9eaBo6bV9Jgv3ybtmQfOTjDrTpdQEDFWaRrn4w/ZAv+zjTmSEN+R47xzgnNSJvp6XvkZP2kA6lSA
35LNyffamEiCsSUQE7PBNP12PkFXn1NtdZBO/6cShCk4payKPSTL+0g4CUwUX7uzF9IjduvopPgx
c8A1yw8nQeEu9YSyNzlzvOUiMSEVz+mtjWLOlJj0wEO5gcjxL0zYbKWUVaGQGWWuInGf0AgXS2U9
07fQ6P1nZNmQuvhI2qD8ZNbw9Ka6pWxovhH0bfyNLB6uXOn/3LB64fRBHfYGYwHcj5L4/l8mIPRx
B3wArkzpdTL4cYIB6PdFW6VB2IF+Yia2nl9iPzOvD8jjmfPWbA/YRoZzZzd5z8ZkxEpMtcLazsPK
lLJ22ZN2tu1GxJ+JYqW0iCfv5nUmTSZpIAZzycNcDodWb3i9cnq94r3R0/dK2LIFp0bHi/1A6946
tAj6rt6uZeVoj1Yi3gJxjFDzexzejAb3E/+C8k65d+NClp10HaZs3CxJ67ggKQTKhTje/qO/q8b7
+Ucw7ZXm7QvL45BoImZVpw71QsXuoQkBxaKlLu4f2Ka2AdTbRBIcrTOJE5pOD6avp1iA9YycaJ1U
+3osgoRftF1TYCopyvcKMluLKw1OoRpSpay7X4/Ho8TtyhrGLjLUp5hJIedZ+vhCze6XnVgt3uYC
5mtlVJJD/BPcW98jt2PutBsfol1zMLfwvSI4WZPKOidWg79LdMn0gK4TiKYtnb5dNaBWHa2I58pD
CSYNkN7Mw3o2ZS9l2YWB51wEd6PtNruEq6UmUQUrcetM4k6GHgBYqndcpeARDDYy/gU4oX4YXNrR
V36s+mMAqJmOMdAyxvX3s3wl3F6zMp4YqalhMfwUsr/dYBdN4LwaO+FvDB00T6R1dbEfK/gRonWS
JjIdcv9xuJp+GeBp/YKzLsnQ0whxG+/aIPUE4EwYi9xH2leEtofXPmbG9PN83aXxgJF0070HaK+E
1ogMT1J+8dNWQmG+117WpT5vEK1+PLvsXARCSaUi7osWMfZ6kIjDalt1tF+6PUQ5Hojs8hAoRs40
naMklP+UDgvlSGdkDJEiLGb8+NVEAUaXz2iMCm0k731Rpoy7iXYcTk4OWHTb0L9qpw7velVkuq70
NDETDxHMnmc8JNs35DurxsLUrCmqvu+q1ZH/dudjCq+SQ66LRpt77I1T+sT2tcfQjaj9UOEMC97n
xHYA8/SgYBUfZhrCFXIkp9ZbxkmlbduHWUvxDnV0xKL52Z996eHfkHN1yYwoLm1mFcapzoZGFXWB
Sr1xCvf9cbpM/ZgajAPm1nkhjxMyr+8I77VTnkzw5NEQ+ZabqDF2S9dzc8+b6LailUNz7k7gKX0w
yPFDDrUCDWcNE+Aaia+vbeGxUak6DSRPnf8xlMa2jvLHP4ImLSWobZcdjH7pS3RqxV+Mtv5llATI
e5MCX8zpv638bcVJ33/8YV2Hb62JX4CnlCb9HMjHo3lJ4dcR//i5ioSFgdAoKDao268W1u+e8PnE
pPM8ja1IIfqSl8hyEiacaVZUzggSsp69/nVL8aXUXl/7cOq8frogh3+hnXI1meFKB1CxxOaIged2
TK3yEDWfYbxzGuijt8z/ixKrsUjG9mnWanUzjjZ8v7gwTfgP6c03rNnMTCn2oHRx9yBo0FCFFZgS
PM/aDCf4KqhXAfWM/Q311sKyPcPNHWpjwQgk2zvzJLcRFnhxkp52yZhtqIvPd6ZJ97NG5Cb59vDj
kXXsFBzG/MvCCrKzVUu4W57cDnoEVSLlR5xBgRGPgJYp9b+4a4wUALJ8/eAsIf8nG7NoMnqi2edo
uv4qOFsg4ox3UucBUmQuBhINhphwmJwk1PkH/4oGHHYPwvkTp0zhDXEqwQ7yT3C1hfXtzJha+VAc
LcbB4XfAzwUib39lhiuMpEbu3cr6Gl+ltMVjpemkb+/w/rtydIDIFuucHV3TzUp5UEbf6FK4HN6D
4tTGuOGIscUHCzKQSyPm42ldVkTqoM7+a4NvP5FXJuTxK2xm9Y+RBR93LQjaM2D+XJYf5N5itvhO
lurMg9V3crKmkH/1rYRN6MfELmlmiqDYumCl0pkJmRrEchrLrNru9uJHBhZfLZ1aX+dDFT2fMK7l
vCSnOpVEmQBCAQ/1nQPZ3RT4DI8iBNZJ+I1xkwOPk+xcTj1w8hfkumc9BZqNeqT0x5608s2txQol
7g85tupapNnpPsT2FFacwkqPd30XH9k6mUnSQXrKa2l86ZHEIY+YpoOi+7eLPn2/DpI1qqZ3HOL6
mg2+3ZFbxIh2nBkV9XAhVKRccrdf0MahcXdH+qbQ22uV93rugvetxEiBeE8BkLbncUFZGMkwOyot
mp+LMmNf+ZR7KJtfTHhgs8zZR9gs4vvI18ec6OozT455xobjJKrJT6d/uyKmnmyqepGEXi0gZLjG
bjzhShrL1PnGeJUQK9HSH7h/n+y8mPFGr/yEh4pP0LDMRLOY9y8RgNTk9GwTZ+U2uNgBCbFHk1tW
rgEkjGoqdZEOsMPfkIMEvCW3NtqnHhRi5ObLygB6n7uq4hA2LZxVkjCeD70clcjeShIlg1fluObM
IDHQE9JT3qxG5d3+x32idC5vjjXw8+zKeweTAAEZv0j0bD+WOKfoKATGQFEH4PUmzuUmTLLX1/Mx
sPXRVkGj5jKEXFEXBGr3J8mdvCA9KOajuseiRGl7cBRBjVpTAWsPhkky2TZR/7UHCuuNAWTy1i9L
sY9Iv0RYc8P+6jBgcU86PO7Dll+ZHhSiPRAep1NV2ZtYvPfwZszMp+YaygkE4hfrbHCnlekYaoYn
Y1bbB3Bho1gUbHIZb+H031tie1ikgd4j7Rlm6KsZ9RbTWyAWPZV1Z2Iwuqk+4MKalj/ZEwDnOn47
yDMgild8EMNQFym4CIYm4l4gdZjbLxHYDSXsM6efx7puDy65TvzPe/FTuHCyT7P6WY08MZDvlXq9
ty7tY7vH4/j1foorCUgslXznKwW0jeGsweczDvGewFOfuKieHAqBHy/dUhXpU1vo7ZJDl4QKuX6g
3aD0Z3rtM56mVBX1jc5kSIJtMHqk6/rkgLrqv4/5c9XL0D6FphpKG41prip3kgcpMI1stSPAwYdj
WAs4Y1Jl286VD0ZcKixNh8pgd6EoqkJkY4jHF+G6AFwIYFFyLcU4hAy9DeaUX3f3uWWjRUvnCtZi
v+12EokjxUSAKxc20xPTenbtRnily9YfpayMkfcpesIcJWLuEm1It2R5zzQLvQ4dp3sbMKl+PnOh
AU1oZj4rfhnlCYttR7vKyCUtR0LdQ0K5xbJs4EcAksoAs+Cbay044EZtM+jtjVlHPIqQiFb3GZj9
yKMarEaCEhm+eRt0UK0oEwrSaTETyD0WykKrbHcd/N6dSyBG1hs52BmLWl8E3SLdFJPmN657etzl
RiMuFmKW4keZ6wQatZkTxl7Ziza3yi5cnz+w595XcB9tM4RvMjZ+FQRsE1MoJdSEVloFg8sxNSVd
Hlc9F/MSR0+Fht+Zmb31Kah77e3ZMy6zhR+GoutuXkxBbBcbbQ2y4FSbfILgz7RmJPSEz6XNXjX/
mroUDeq0WqTrWM50V7GBpVtHXl5K8xgTL5/gERYzJTC1PDMuSWYDvatAOgBkjPNNpcQTKHysXjwI
R6dbKqTGINVosSxVC0YTrsNDvdeNesiFeA5JweMNYOr4iGQLm+u9Sj+qhwJlXhX7YxVQGR0lHE2O
c+g3dQEbCegHw+BIW9TpZ/XH1vR9oLMr+XvFbSHCFc98Vfzd2q67UuReP8Vrh220PxZt6I7BTVk4
KGMqu07CgtakdTSgsdNuTkJEkpibXMmgA2GXChE19ce3RAxeDRLw2ZtpngQGUKC6l8VxgEIM6Hnb
XtDVbyX7KcgaqpXA+8SM7UiY0wk3norRhFVlnaTMBZf1bzPpkIKCqvkr52q72or2fm4DCwRkEpch
NPcOOLCfl1y5AcExMwSRts/qYN5Dni5EFGZcM4SQfXjUcAfpnABX87/VJIK92c0bSBPai1ZpJ2KL
QDy6Z2l0Joqw7DwQ5Gg8FdNXYx+ALwVCCj6ALDSsQTlhWhzpKh3SeWWG7lKmaq1FMXwVbGaAZPDf
+CH1BGeMyjDBw17EUYDecBEbMaTYrzS46OA8SO3hL2wqU9e67o0V5QAiawCfbOBTRhfdPLJXFFMv
aDN4OHc6IexMI9u8ttAsgNAxnMzvf8Wjy2LMknSYD3s1lv0zFCZNvMHYuXv/U/jQcHpNdSjXP3c0
ZKTJBC+GiVie/o1Km67bsUPJAzerpE6ZONM0xWosJK0nkx1siMBOih6cA0Yp3ywBFZzYDtXUnnbM
WpAT7ZaNe8inMXJ4Qg0bO9A6b0NjfrodAPi4mKr0E3nkFv3tPvgjHhlk1QrSZTI/10zcRuqh4K+G
lpyw9bOH9g1XNbgkGCDmPZX7LQkVuSthcfQoBTFGZjbwDEWUW3nGCDWD+SUEY5rcpSQP8vj8xcai
XIq8A4mhtnfHkzncyR9HutNdpzFtkeOO+qPYhIjCHvwlJPi1LiZ2MxSU4nb6yWlKyAdhBgU9mzjj
jn6VIhBou+EN712nd0M71NU+CBq+2EIh77bBewjg6FraMvo+BT8iHo7bK4vml0uXiqmJ3H2P/GOQ
D6iKjeLtz6xcGqf8yaWVHMANCcUF2c8DSlcPpfvbdIRA8YSFtIzfmQdafhn47oFyjY+EoNjjwzfd
+QRL3y7WfY1nuH0M6ptUI0t7FcLtMHs9OVEokbcblcKwyoAiEepTYe0NviyLNTibBd+zBrtuLBaL
H+0bcrrMaeKNhZ4S/y6s4Y17/bmqdp6C4GAohTsDaxuIWOHhr3/FZFOWRyEU5/wTcTTpiDPuXbKA
GGmWh2Qbp8zD6qu3bXa98T5pwyJlD8U0nYCHBNTuBAAuNlUYiaZ+jnh1K3qsJCg7q3UxNJu7pGMa
tTqQxj+Vf1DcqH0KI4U9PsxLnZLKsGg6eK68kw+BiO0bLqUtkKp0Of/7vVISS+uZuoVkccKjYVMj
DRr7QX2cXcKTB57e+iAMjixv+BdMuo9H5arVkdvkdzGDHPHe9By3xQJmbJ/hDay4evXGOgqJvpOu
YsCvkHPaJ4kuhCCE7+n0I1tR/RD7JfDEMhFlZ2DaTXkFoiko4b+5psdBGXAlGAPiDhU5vC0C/Ozt
S1I/JzAyCLVEVw4jMuCO5cY4Dlo4N8vD4ggMFa4cZHzfZd7ELJTLj3Wvmg/2emrl4QksgMdNCSE3
eUbtTkahXm2u9i0v7nC4AmKfigt2vNCd44Mtc3a1T4ZlQeUzMor++5RwZCqvo2BZo/LIqtvoQWbT
30uenQeA5md4iZthk1oWFIf4H3sLdhYNGRjBtNQkQz6G/sgjP9SYqL3Z6i3EMDVM3tOUv/QiqLNx
pi4WmSTVBrnRJa6wKmnavipdGNdriCUh0xlTUY6BqWFD+dOcokMoCfVNnP6fCarZ7Oi6wnoJRQ0N
eaxb1pCQ+z7JxXpxST13TsKiPp/xYAGdvkKz/YUAgLWSN0RY3UrmuDLE5hZhXctCZ8XMmyCBwc79
dxq8gbXjD+ie/Q3G7p4WFhHZWse7Rp7RvUJd8QD6opdZfiPvsPsOgFsGXg/qcN6fATzTJDLQJ4rF
SrFhj+O1FIRWZ9i2bMisOR293B7D5n0vO1hIpnlPX5fc/E30VDAPeF8UXsBSFotUSEB9uElQaQiC
jXK5kc9oymFsP6LehfCVugtIyCxnu0xeFHoUbDi5tkO3bvyQnkVCbFrPZdMxqRC6BLHhFZsrBj7H
BCO3N/KzSZv28oiuXPxI7LttsHCbbXDXDgA8+gkf93qU0DTQL5zu5m0eNZch/298V8FtJxxtC1ds
Sp5PL1cbOCHZZtw0ZwTj8IWfhdEhE1kzsI6XQYARbR0kf2cOI14jRjayIpkokdTawycFlZ1ojK1M
9tFOg21w8C0IRiRAgdn5F4ct3qgIRd80bV+EWEBI/2Ikhx7mZAvjsrXwDvowEArMvTT65VvpkEJ1
ERAcwrAW7L3DmEkZhemED4JoiJewyVjAJq422tEksBuCm8S75o0Jd3+9ElE5zhw/Q0YKtB21BBkK
o30mSwttYzPhetlsB5ysH3frHp4iMGHbQdhS/kWqfTT2Hbn15r+w+nKE/Ggfo+OlA03N+KF+YtnO
9vt8todZ9LqnDq4OobBK3HgfcRQOjNIA7/iZAIG3VWqJiVnabIqQ3HfO8WaFmem1Sac/XzQ6qOhR
4cm+3riCYTu2zUSGz7D1aqC+voDChJ1NeoW2q3MzMiha1+0vXVtNvi6tr0FNM9lrQwRONccykWSr
HlgPbhEaYnL+LVZCmx15pleWix+higrcQgTQHc5UNxc8w4tUcQWgcZme3eAwlQsk8Xq+LIly28DP
dEugEQ2Gwb07E8azuafxepX2bmKCseeSHyIQtUMTL5jy2bwDwPLj53mXdL0ozSbR8A3wPTqU6QQM
NJRf+sPaWRI/oi9Qnhgq0Bfj6K9DIGQzTuSqLuT8pz4CED1RRlwtElm6xzUlONIqC9MJ1n4glChY
8Z2zfe7YmsPtRXmQ9qDcqubqCEVID20wzIRPQMdlYAl2X0bAkU2lTdQXJOGx6k+aPY+rB4aU0YRK
/EXcW/1fxNk2EV3oYz336FXymRuDMOILcZOM3bjLX79pJ1gSCpaiOzaX1AG2Lj3+GpYqGjiJsxg8
KzQMyY2dFGe3dPdVWFPlSrFH3QvWKh9ijR3cLWiJBDArWolYfhcQCvljKTWXg3QC6h4zesRgr+In
pdbV04Otg3vHpWPuAEX7D8uOsxSyg+0Cqj06hHQ7DK8zkQaFjBFoHgzKpu7GzkwRhhsnxVUxqLCZ
SCaaIW6c1uh3XU56P10RQbO5ci2JdAWWRseJn5NhKWJHwttpGE6uqBWgOMVu8i43lp7NZbYbdNbV
ylxNgBYZsDrwlao3Vg3JGjBfQa8fl7ecFA8MVRZwhl7uteW4o+oKq4glakYXW9LI2oKiNqc39g7W
dm1lytC+seCQKStLltuiXZs5fWoLohFY1uk64Dgwb0MXrHsGI6EYjBVHrZmvxM0VywsCUoX1anmC
nRM9DDcLaiLo10xwKnZJtsyOzwBkQ4hrRjYkoCqtOgY+QiOnIU73BDB+yTEinv5z+2AMIUnFdhN5
i1XrJmlH52vDU1ClvKiptDLXdb79zjFkhTy56CvzEo3F6mcPHUuiZIw0na15xTin230WuRn4OMrQ
XoYLw4Q0p702JBUDtrndD8gJHZdb1NfP9ycDqzrKXk4829qWGJkRIWWVzDaA3B9U0BYxga7L5kFZ
+o56N5EvWNIzk7eD7MblyfGxMaFv+EfkzTuZ7jJX7trcvKeW1L/mcnEyD0cVJJBDFB+IxVtXRZlH
eZKVLRLmjC6YQJLRnxxkoJhagJ88G7bnLFXKwTA/mhAXFzdG2E4LAVj/ZN5m6kCBUMz4pPpasw+P
9Ggi/w0IjocvZtt4gQd6+Icoo/pa50dbvhaldAXRBZaWoTtV63lG7YW6tuB1w6BOkObz5uiuS797
v38wccwFsG2ecLujkT7C+0JgxdaE1dJExczoJTjBkPN0XiFF0Cp/ovwZ0pAtu8Nz0rC7JKM3Fej4
duTO7JLUXFpft4sPpiggCX//SLO74XtvwIzP4yBxGwPIegQKklhloQkFuE6gCUH4ReTq0fKHCYth
1goUhxWeTF2w5XxMvdTMXutmq+oBQ3WWsvFdIS53zOKk9/yfA1/PIW1g+iPPhxCkRnPxwOKS7nOG
WQ40Pvw6lw6HZ6rRiqEFC+lRUNri8PqKIGRDe+hVJB62eN6VPo8itAWOOEB4J15bv59Z8TXVajMD
DopdZyLuvKz7B/fVDNs50rn3WxeHvmXQcVQKACPXWm8bp6s+VONZUjY2Qf3sjRUcYSiQUl0T0Uw8
geVdiK22PjPLFXODsgL/hAED98O2dHSO5jTj/ivdEx9+gShJMp/EFMyxdlIedWnTzoT+z3xWWdN2
cNodoZBITc0e3vRxMNww40lGiaQ0kIi0h9EAUp8J3pF2nG8R9SK5avgRdR8YIgFl64ePUf2Y9fyn
xUPUqLVhnXrqySNS8cggmqgR9wLQmmFOg2U90i647cHKoeuWOdAll3byvSbFb6RXRbNp27f5Ga06
EDQPNNx+7nvAGS6f+SZTFvFzYZuSKNzDqAG8UgKr5tUOxU/TM2shd4s3s5LGBXpuzi0/wX1VBmsq
oFHBKMoY1qIuZ9GeAnHNy84eJIj1+pyXxqi7p3TSxFHXe2xxY0XG9MFenRE0+qxJUHPbp5BSc/gS
9v+5UfsBq/bEjxgx0Km5g5eNh4nr5bBhvk3AdDOFzNOlOHsHS59GUqLj0ac18jZ8nmqTPTne88uJ
2dBF9raTOA6jxUFjKXzAfZ/dy9RkSKus7RDrXKSd8q61ru8Lyzf79CHSKBm5QqbZ4y/dfI/QWTIC
wDkn28C7i76dQAUCzQfLwLep/8U0WobJvkvemuqyBkoNy7hkI8kz8sSvmGjCL1BG8XngVncw981w
lo+YhWjILsplOudTvMeLhhtYfoL8ROf6puLymr8JTHYfpvEW7mwyCqb4MmXOKHUm6SJFu0K18th9
9C8taN4LM0pFhNSjks8kGnjF9eyfofy0i3aeImSl9ZOJYKZWawp4sGQvAyR6qmASihQCMOrf6nin
JLMmidAXxI4H8iWdJNqOr2fwLTYjAJXSWgfUMdUD6mtDUp2mxjFbuNnz4hkBM9F0oVLSX0hRuLdT
B8lTClrvG4wDcVUAyy9NMMxZRl5pv0aOjjS3T99f1uKoT8MbUnj9dKNKBzmtZprZAyR3Rx2D6lSt
oMrbPezoQdqZYpaXjSzorM0BjtrnG/rah+XVdYdJIKXvYjw5VE5hQqzU5UiTPdQCivsS0D/SdLeV
32fWuLcxHazGJMwEppvVRhI0XSnMPv262D5kDArXOogqTnhBkeAaAOH359VnUB7wj1Zv7CWP2zmR
Uzqu26wKlRb+gAZ2LfRiISXF53nG85cj2bELOSxYyAxKLEfPQb2EDpiB+iwSzbS469+Rj7bOENqb
BpaJ++B6bOfoBPYsGLCtbaw4/J4AXggX2jhnJG2Uz9xrzQCRjm+BQKMQYIxOqzp68iKD439bfuyj
UPuN3U4Wcay+aXWjoWmyQICj1zUJfnFmCOpeXHi2uoaZJkGF35Tsl6YQ0cPQjONJ4NyfcagFHyba
37GBbMHLkAkR8QIzk87lIxQQNtysMWI+YnoyO1r8/veybR27clQrCAXko0SUrv5cO1VfMFklZ5uV
PWBWdInvRg8yFhGVhwVPo/wIs15AS5BBRbZVAyJDWvmQSB/mG3YtmhB+f1g2XDunYPxBghFutIxd
4eKEO+tSmWBU5zN0lxJALCVD2OWY4TKqjcJbyNFwQpmTWabDL9gOn6zLCQCGo2s3hP4GQSCRB8VX
d2N4Gz/42dsprlqJ3z39xC6RZiLIZlR6lYMd0WRrN2lObz3qpgEW0We0mg7khsBZE9xn7jA8HLFE
6J/URkjwlY4PJjBCm9xblpzS8t4qxc2yxP1m0kxr+K6tebo2D0B9ynfOvGscUEc2EN+KqOnQ1Wqu
j7vYB1fOoGA6p7TeegIf4fwl5HnHL8xXQlyyiLxC+wcha+ZiefTiK4yESsgnHSWJ8ZuJHszIaaEv
JrqTP/7ry+ZHRw4mpnpjdtsJFpLzAVBRUW3Sp2787yunUjsx/h+S+hK1Nz6NEjdJ2PXvQM4OwYic
t+BaF0xn56sQF6Szz3vabPL+9JWu2AYY/7veVq8/4EuFdGexz6pyYCA4B7/qAMyGllfuQs7Io7Jm
RGNr7+B/ZnFYFNusrytNVCOhZ7AvutUv2+QJr7as5irbSitEXEpWhp3iYHQ/B0IA76TdXYMb+srH
46bx29t8kfzZUBIbq39+VpU/RKuPSqw+GhNto6phgUuO3qdlr6c+MVcfGgJAQYSPnw2RC1NuKXBR
xRTMRuEKtHf9dYPlCVrBq5l43POZuOpbt7sYBZ5Z13wFXtdcWPaapnEx6l4jc0fWD1egRx2VcEGY
d+85YzpZna1g3FlYXLg8612mbpvZiCSwPGjBQxtG/QURdFPTHnv1pNXsxzHa3516VlyBimxmHvTL
4/HcZJqfAz6nVCKoAyykZzIAjuxzlXyC/WjAZVQQSvGRxSkhR23VYVU1rGENdz0NspYjAMM9D3fF
Mii06BjUChnrdo+bkdCDHndj0d3IGGSqV02v+wwbMkYHssVUfBtjQV6WznLGBNLqRPn3xcqj2qn8
2SL3Kcjy94VYRamcU3R8WeS7VaMAJe0D59+HsMimkY15qQy7c34L7v6SAR58skc7gi3khV3M1lwO
EGUVJekTY88IZVZ2F8VcDiQo0DeiSBDNNUOzAyNB2WnALAaXuekcsuyeZ1uYwunuuXdsn2fb9JDT
K6JRDvX9MGIdmVB3BPNnHCYMg17PHMTjCLmd8Vx4yrJZYnfyR3s4O1Rw/DBZ980/rBaOXiYNSPoF
pkEijJqxi7e9KkhebbC7gkZ+Cpqak+RXUM0tP03jvvxFP/W7yfpjIp+1Djmkk3LIieo32ZFWQ6tF
RgyHCItqer0XV5bWj/I5lmSy4HnOrv9HdSjdBbWmElv8NStBtzJ+/l1M6q8XMYUvG2GUXvHWP5Wq
DfqOXfXwg0aWLTXScRFT8U/Xg/9MQBLO6cHrP2dZYvL6DjnoHgwFfyLMGK+IzvPl2bmFvA6aZFqp
+i9k4BslQG6egoARPMIbSel/ETqXwRY5YrjJFqU9RMhV09AbbQ1V5GtYWhHphNvHYdateX0OFfu4
xofYU9A6tjamGWRphUlLZJir4pIxvn8C1bOa5hQdHBJMsU+GwL6+aNovDcNM1s0WiUQNqwW+q35e
1MNPRbCNQXwFTDoEYRe6DfbB0lTM1KUsT43WELkkHth9N+v9hqhDQpbBLfgQPLu3oGgyMTCx1N3L
9HaKC2nGTA4NHuibYqvi1CZHbJ8pz1E3pzzFKj5MgF+ugjWHf0HykGtkKhdvLPRGOMWlzQFyxhQQ
Ot0Acew2+qXKFkRaqcs9Wg1z+wtM7xOjA5zcpfduMQmbmk4lkLm/NZWT3EOj5pOADlK6/lduLAHL
xJaonBPtvoVrm8M2I4BZUvN4SHWoog4GQ579klYg737vfeJ/wQu1lB7AV507lLSGjZwm9raCGrE5
CX/ZiQsmymHTkgd4mv2ASYHiu7N70fzjEOXDqMf6odHbNetTEyA1w+OKKdiGg6So8ETbiWBJJNpV
K8gPSi3c4762m8BY2HAvgEUe5tRgt19wTLljLwh5WXV2OSE3C+H57kyr3ox0dEiDbASD3QPOGhhE
0utegcUp5BNf+1l80z5zI6RJCi7Mi1yP2mhoOU4S5l/CZTaxVIbQt0Vm/NjAytL/sEYGjC263u+8
hsVrC9QGOKEWSskG9saQrkdt3TG4DmGLso/7r02yTpHo7U8xrjuQ/J8P4mkbZHwgVjLX28UcTtc0
Ajuk7VlexzIO4cY++tvxSxtUyPJM2YtJx+GXqWj/9bp6GO+9BhOSjF325vs40T7Ld+52aiM1OAdI
n4cXCkvTvGMX8Uvzh7PRRbZTIha5Zceb9Cgx0ZA2VeifO5N1YNE4I6sW0/9V/0QY8NSccMUOPZYD
0b/qIsp43yGQZxQOBKlCH26aVOJoNQcBqx7u0SoqSGhirfOpIQImRvc1pgMyOjHSJGL6uLH5LUI8
JgtZGV0MR1Fg9f6N/vZWRzvoW1PAiW1SnqTX2IjXAyUydsmNH9g1t9r32Qysbzkg0Qv9fO2q4vjR
BVtPRmZbtTBQWMnRSBrk0aRktF2Sm0i4V3+INPvle9fMlWqwsdjeN09r7wl346/bVGbyfDwVnMhn
dOOT4KlnzXaoAyB/l21L40vbZrd6TZuiuk4h8BH9u5VxaG3s4SB9pJS5WOF/vSj+PMYeW6M0/Hhl
RYb8kOR1dRz8JaH7nTxER3sWTi4YvwqMtJ+u4efuFkdSf1CxzJvAsryJqlsjngH6Fif5I5gXH2gA
pGFX21vpBFfwuY7LGliKWPu8+4/7BEkEzyTrcaTjGhq9/Na7ksuSupfiHmhnY8Ch5b9qiMqfgTtu
RlZSMfvn4scd60LwnnQEOymbKz14d6UsSXJSz53q+Z7w2KZUqHfgE69BRgFZMhamhDTR03Z0txWE
cN/Ayg4zTebLequV+fsROceg5z4IB+DaOfLn7xvSPlrV8muLe+iE2XNgS9YUG5QgvaT6z2C9rjUB
MKUR/YUkA6TnXS1ko4g8kZv5UI2y3JlbgN4BOUm2MoLrFJgJ85jZ/HeQRn15uWPcbcEfqfUQrfIa
Ba3yoXZUNpd8IwBSBCGHbFxnbbk1y1kEbvo7oDZE+W+QlFGECep9EUPSmif4JtzeCsiXhFJOBkNG
K3FWb/bT1/Rd49wS6FDdCIG1JW4y5/XhRqgvHuzgi6PsQR78U+o6Td9E6cfIwuRfJp7YkgD7+Azs
CKiprwQq4cV+w+ygY5oJM5zxIyJBidMtur+lCa2B28hVIGgG35IYYlgMdF51RNroDI+fY9FkbWci
XAbsp8flk20tE+EM91/WF8H7dH29l9xZWerrFSc33CryaxU/sCrtl+krq3LTo+KAntPV00tEglPC
yur4ZIYEswdr1e56lnndBXhlQGzdsgq5NFMVhkM0KZcxt6ydRyRcVOVRK6HYG2JcHfRcOS2eSkc8
fAeatjhxUh5r4yr3I7InAtBEkv2x9rUTCkxPxXcewauBSxBQiiTnsQDCU4uigdS7Me4S8FdCUpbN
8JsfDEv9rTlZIEjxQ4rkxEPLGuNwAEYdsqjJ4UtA5qlt8iExnLHVndBvT25yeLqIuMxbtGob5PhZ
uV+M0PaTwdCdeZl+hHShh1yMXkev3mlmLIHFYkwciqe2goLP23o6INLtbn3hvv5RzlCghYTo4yzt
hJ2809I8MhJYwGGLLcSxTu7bNzN62VkX4BmQ3FYt1K5AfMJiQaKnQIGzLusxIxyAvWCHXWYNHL1d
ZBweLTnTX90Up1Jh5haJfWGUO4WT0M2/bYYGx7Xqh1TI4RssYztySPF9Qa0gVgyQbg58tgcrrqoS
P3uodYJmlrnjLqxrJN72OD7DFv6rMRN/Vkchx4ty8Z189Q218IdwwIqdD9LWuuFW3aOIN2MW6Mdn
vtdNBslgb1nr0u/hXFtJIAYTkQdu4LuAUtNIJCNbFbRPQKkgLwLUq0WGBD6CLDNVLTxngesfZTU3
fMHHUnDcHtGFy4c/ecDq9IO1Aj/V96wDTYHPyJTjPewBAJartAk0P1PzI7V7iDno05sdkrPCs0yN
go/3pEDavowsnR+8WSSBM4NVw4DJ0oYrNRcTEs893dmxK8R8cPTIo3hTKeJx5iGT04G2NgB7HliW
VVGH4kVD6F1hVu3/eEEb8AxFD2YEIbuErt+NmEbLtA+b8VmATe8j6i7fm+ghAiz+QgqmOeZJuMMi
1IYz9fJ/gFpibvXtnSts2F4xHiiGIw6uhRZ4dOFdik2bS8jFMWnaf7dVFfiR+QB1M3+Q9ckOd898
WVr1EIgW8bEBheWU2ItCJfUZLlZl4HsdOKDw2O68Cp4zIlZVfHNb/ECjrxAiWglr6YA4FgAJVGFB
rMhuKdjl2fXSsfUzFTkzEcRaXXpTHOWBCbefdHPSy3jx/bY4N7utJpj4g9uH0ucUqlEL1mL6PRPQ
mNLmzDgr2BKK7fGNWbvTuIhR/KaGmLl44rliccPVHLONiAik6pdUjfNhOnhuJ/sROm6p+I5Jzg/E
IGc/xnKGovx/mHUJ6RNa7R/0Ec7R1R3l0Rz+/1sDUeT4+uvuSf2MIZB5hwV1nMhMEhqPyNLLTKYV
AIlBXb918B+sG8NPzy6tr8KaIpnsJmc23RFLLJx4uqaB2QGqSi1LWfj7k+5x5G9PYK9bSCNDsJLJ
NPfShpvVOAfclwtY5PR/sWly5ci21O/6i+3rR1IZtIspEUdCRNGZEyCI0sxW+lk3G0vwGLI+OVie
Gt/Ic93v7EEsniLsOdXfbGWK/w6t00JhuZoPAxvIHW9hjq22RUadsGW/5OOCw8Cjd/JKHJxSSiWK
zcSimOaWVU2Sl54g4DOMawvmeC22wv0lSk3dCpzuzB6EsWubQnf+595dMkpg5bfd6xTRCEAw3S9d
GJLaZjKbJpXC0HWrzFATEQmsnIwcVkI5Wc+Saoadnz8nah+3oSShd52Rq3gWXLIXi0V73DJJupis
wKsPQUWC88hJ3psp5iydwtU1qv7JwikIBYyUhVwQXyFLsFct7gMmpXtu7fRHfzaxqFJhSgQn3h+A
1lfIbKjpHXytWH1BRSVF575Nl2xzeXVkqBN/o3gamed9Lv+8zVTRtT0DS4C3gpKq3z0dOFvmR91E
lNPx85JOPREMk5okJ2Esc9Fjn/U0tqemL5jXN80vnVEG0ibztAETF+v1pZbpRhZpTksU1ifKx8VZ
ADda0soYR6m7qqn5zTJzHWpYEFuLChc5QScUSo4r8LbH5h4c3+H1A3oorteFHqBWVajpIDi8842k
Lyg9XIoRCacOljrpU0tAtCyYI/+MWeCA0Mgf51h7Ff56+UHpe+ubHKFNM8c8a6E2oiHIWJTM1yaA
jfcPGvHA+2kYMowd9MOAo86XVyYOIqhbXL3ERWrYT7mKJ83U3WJGWngtBsFXphgmDfmZp4/OGjKz
OMs7t/X8s5y39m8LSZxi9w4RiNoroBM67UtyauFbPt8s7A0tKMBkcVGOrkO+x2IRf1562vz7sUop
N8HqRDKvBVQuYZ6Mys5qEuSMJrb8B7/EL1XjsYXIb9vVgVgCXvEBOoItfHNiB6zKe1eL7G/+9RXy
ytcRvMXoPznuZmT+WOceTN9ggRRMgIttYLGlwYwJR6sKMsiiqPDMtie8upG7LY9C83UE73BaBe30
szD4CEt2sZiQwF1IziFBeizc7a+A5apJQLH5jmCkgnT+6mWbProC8BIc9tWCHfPXSfvEfnXnNboM
CTqmGhMuNeHbpenv8QJO7nXrDXUNfOSIKn7opdvShcS2TCmghRP9mXSM9dgj8D0JeTSghXrX51wr
WudXoOa65ZSv3IJCqTu7zSNWVcH+He7Di63NYKvHFQXZqMvIOxSik8nTEU7RNfIfvFQ7RX4ytRNZ
NJehv1vI4fSgYIzBkobin8MYDm1F0vNEQMtmSfJS74l7BpvUpSp9LfqVNABU6NiesnE6v3sIdgFO
17mi/wF73RCz/CC2RI5PtU2jHg+B4+A99k6POyDASQ2aKK0rsV5Hmgpd2fcG7ZZo+GCqaZOUson8
t42ENiLE4FZ0cOCn9WhRN3DHO7mbbmwcdyQQG3Y1ZyWEAv0QVEsoWZghIVadeKcPs+qO/iBrah2y
IxtDBzs5r3UupZurutcEql/zlBKK9/Nyh1c6a/0fcpcdDoyypVe8qHoMw3M/7IoRwsveqz9a0tvu
w6OIhC6Q/RP23SnGJNU9P59KQK2UYXZ7wr263JacSYWMlmCZfYX2Mhv5kiFRy11/IyUA8rJRpmtN
uxI2AmWfS8YDdpdJPp8hZWyl3bd7QIPpVHf/9QUp4ufLD0vYLaf1TIkZ48qc0fimJ/2GPkFdNDzJ
QdTxTV7/jnStFfY11jYSbacguYEZjfQ46rvJu5uAQJgh5OtwAfbMHRLSxLzRQJoMbD/pDJW+0/cw
9kBWlkvCW8ay+Fi0ceIOcGC8yicAam6ai1iwyY+3SFCFoJuuxgZi/Qu/cedpO2Pvf6NFJUeOL/iI
OTVEoR9DPKGp4orGVWjXwASOUbTIRnKJ1raNTTY5GL667fvZBI9oe/YluYQ2FfRHNcQzQrhOxfg9
bK9C8iQT9DNgpbkZAglG9pVZshSq6j85Tu2hl63uk8Z8OH4V+uzDLDr3A1bG6cRRwmG19Qa2RsLg
5uyw8AxdFIKYDgfxr5iAvtp0jUyJIHAo1J5brZ4zZLG3XZC/LzLgSdnNiWGn3u3beej4IiiumOoY
wt0ANimxZLeyo9UXf4ZuAN44ux4uC+R3pK+liPqfCKVqDH/gevKO6KrMwZrvRcNEyUuce+/2m8dA
WBccZYSbl9MakJdN1t1/s9R2/G8p/OE3aVcso+mgmSSU4YC5asAlAbifHpydjAuVUHZvMyWMCJn2
b6BkU4T0tYuEGMh+tJbpOYvjvYPL2BM2prb9y+mhkIwWH3BKvKzjbT+Gx7MsYCHd5KzX4P07I+SR
KCXhap4Yw1pq8JR1OV4gqL6WWujbTYK+pNDts9TjKC5aE/v87ICQN07DT3TpzTEf9iGOOesIuU8m
bIzcbbT0hESnGlGkuVsXsPcmYmwax5WyTomI9sjuFGsfGWTlQZUf0yNq9sC+ii0biqu5aH4EMGx+
zLogP5spIkHlBTOfgqB59qCkjRCgFejlYM7lcIYr3BdhGzn9E/Z68M3aEVZdl0FxnLvO72pZki5a
UgyQMxIJygBW+PUKO+4548RdS+vQ8aFedbA/2WA3MqCkv6nbkGS4Y55eH1THszdUwVItvz0Ecdr0
Qhpfa8WAvsuYu429FYyi61pHfsawnjckDkzgrUGczpSPO0IVWAskrJYzRyq2B7AWD6G7p15zTsmj
nEJbJcd8RaIoMYYzCmyXS/dRoUa49OQJvLn3JQJiAOfeJvFrjuYMOPAbI1VFNC4EMfevtTW+0lz7
p+nUO1nbwFt8joitEbKIm3GW9U4Abwf/DV1OxKy0NOGzgJMiqShsTS2/zXAt+8O9E8hwUblde3vT
tBMBbxyN9MQOJ85TEUYNhGwW1D6SB2kXCnqPKErTsENYvqxESYBrpbuCcZB6RWI6PNqhF8J5f+md
limq3Hu+ahHIb6QoP1eizb8pQTCGAdAJYcRTZjZMekRDsQFE32pDDFZeGEzAWDzBZ23R2WUllUnP
N+ipYaKbRdzf/3qrjtVlP/lI4AK+vJpdlszb6OT2NmuvOiwKYTT+viUnxgGLA1UQrw2CdFGHREBj
rbs0SyqA4s9of1JdzziI8xipMcBqNJcOi8YLzC3ULT2i2k+/CRu6I2p9y7NgpGNIY3Plv/W9aY+B
AiQFmFFx5tu2Y/NgOEtNFD7AtPsFq6AhWUSIucjzU9bh/oItPdOzxLfACPD3dxtOF4UIYs9xN4Cd
hpHq5bRpdwUIHT/DUs5rB/MMjeg2LGU3Ppt4MjQdxg15hIgMQ2TatzHFTjsO5zM+FrJusXMD+aDd
63GkofmqkocQCmUdVsUCqhrWG+jHppDVN4N1zyn0I6nS/mxRCwyNP13qmcaG47AoOEtVjxlBHxFN
/9/lW/emxcASzZekNTVSY3U8yP6TL9TvrsFP9H9zAYZZ24/mCSpv+ZxdJHHAmgDywcZoFK0OkgCW
MpzOzJK9aSzSyJXA5l5R/HN+Bqim4Ug2a7CdbRFYwqPT4NS6kSARafIZkCdfUV/pUjUjrCk4YBM/
GTSItSEZ60flbeNnlg5vwwniWA429EK0l2eFBX52azSi9HkWLWZGq81+N7dV6SwD0H9OcMy+Lx5z
NjyOLsGn9EHfFY3CUe99rdYFbm0t+k4tmXkgUpes6tgJfR4zf6BuBYl5SY+MvmRwIsJuOB6OKwdI
QR6Nnk9N3BMDoAH5cdmV6DD6rE+th+uVRfpcsUb1i4vNqAdVPzr3BBtXLmQ6gaJWyqmnti2qoIjY
fgEBgVPsJO1nkJnHa/wwPP4t1t5BwgyXxDIz+ZjkEcRvXOtvMMTFXNLqHfmk2iW4GWOEh8d1xD84
h8aG3VAbYvlRpou4pwNHW2UdaaQ/5FrkoNmS3ZKENND/LUU53E41mF6rlx7TCHozmcd/GBgOM6Jc
nZL+YaRqfYxQdCQkhR2hhf0fNVPo/8YW0UgZbHJuAHEDAIj/UZlpXxg0o3fU8Y90Zr3NPHm3syZV
2XppaKNSCYX2BZFrnpRUlV1W9jbp4cjFnlkNgBRMjXeBn4SpuMBvVF4vHN+l6gy2hMhAE43KaZ3f
eSF6/lakaHQxXLLhrqkWxs+oNOBTsVvoAqph6kCFC1kvsXKTgnPcKotmwDCxxVj4AlDG13eNPN4r
MrxIDpIzgZ84Vvn793PwT4ViwJG2QhB3bHq/3fqHagBOnprue9LTMMRHLPTP6GD5tb9YR8Z0rNQL
UG/ljeKDhBWkcmyrTZ7NdARzUEnVPt/DRJvFnH32MtNAaA3d3BS5De7BbYVe5aRXHPPX6S57A9om
9ycmeuvCZjO0Bjx9juMea0K9cVZIb0LPhIpJCJCwTqxNOKXHfpT0r05hv4WfhAv4m2vvxciD7Iph
s/T3Tz5bKc7/+WN2g+0+Xh2xHgRWDFky7PW5fTaaYX4U/1Z/jsg6xw4494qJIAZ6OOc5kyC/heXe
5Bp6KE9VhdnfLhPMpg1BAdTWypy8Xu9uXB1HpHDxrq3WDwpyrlnYRg1fLsQcI2TpipfRqrcASulu
xj/fVmx4Eudh4PqB4RYYv176UIt1xSAOkySdd7lApk/zhMopDVDjRmrvYgxg7oYwcq5Nuryiap5u
f39WmGFyp7147+50BWX+1oK2gawlNZaawiuaFdrVPoLmxvsM79OxM5xsFrJ50ngwE1PzeEv9zmvW
hfX4e1CtO7lyimd2KDAYLRq9uPe2soGTLSVr4UnyD58+HVUghYEsL/pYJOdafqSD0eBSaTNPB1Sz
Nwm/3fYb7EpVRQnV/sNmWBHX2CLwlWy78O21ebtsYkjmpx0UzDeIuQki4lAIhqCY6E2OJaI+rYtp
DKI2fHFOlmenLLbMzFQdZAg0rnMs9vfrrmlSmwEclqf0hdZpNYUo1EG6bY7wxTBFJ1exI250hK6t
l2YBnc8t/vSmAzwbU9sv7fVVK8SsZ7QgGQxra+jziPx3E+JKSS7rSonFJyfUI2bJ9Le2ycva1vMs
5PrA2nHOa0jOn+70LImmBVyuU6N2MT8SsuBiQ+T5VFkkus72pf2Wo2vXNuOM7qb5MlLzBNFk+BSa
IvYTV8Y3Y93HsFp0ys+dIzU/TXT5KeSRjGoLnrBHivjtbsPk/Y7mgyI5Oog5sWx4GSYU9WO7kXb6
XgUUBeOIG8qAUJCnoeaBK6Zgv/O2mwnomtg8uMDInsIiE0oy/z9PSjlkZk56HH9bC7aLTLi6ItG+
Dq0vGOpFU0noeylgjdAXeVUlXuCTGuxltiw/FKKW+6yrwfitiLvW5WEZpKMz/LVlXgRvzJBHm96j
KIX6hFMCVTJ1RR6ySsJTZIewm4XC3XMtazs7zJau9pAxsbccVCTCsk27y/CF6YreV99XsOnKYSSl
AwboxjSC/qNOTZ+KyO7i5Vo0J5OhoETn4n4q8Fpev9h4N3ZlPznrlp5en9IEs49C0J5S2/dxXYhd
QLLFzArvgkb5V/4if4pcSAoJhAnhGHujn0NhGuHHhZhUb+9/kTqS2cANcku+9wRAfZURMK/lRkdR
3sWEY1LINetoqKtlSRr76VbfvJHzssnUgtSKv9y+ZRYyqR3GHJnva2cKea8Vb4oQUVbsqLhaorvz
W7dAPiwLtIcf0pbnAwJcJTn85qMFQAVWq1hDDL7WNEGLr9T1oXerAXcR1n1JdX7Kz5NqXB1FdjYw
EP1TcuaYbFKSJ/JTVZJ3FqZlVPM74g351HElABRwg2OdHF291e6kqJXh2xcYPAomEVgDNqljjAIG
3wo4+LpLHgFWy+Wdr9PwquXv/TuMGD/4djJpJIidQcmdolxpXKrjvGfAGjXZIrFslk+81RYulkIj
qZdX7c5HfLu+S1G9nZ2g0RoIC+86EN0RG38pNrMoV+z/Yz9axOaRYH0ASgT7vdjzs4Kf02t0SjFA
IoeotCgDORCVLA05J4av27LVk3akSpOvJrXGrJcedNpFtedUvjyO8tByMhG86d9XlxjmqWtGuAdS
Yb8qh5PTe+Ehl7d/bMhkRAq89kz4of2oTM1DkVirPwVsYkcUcsRcWruyOlG4oIgpO5MdwfZyooDc
gn1SXsO/M2QJmq6D+3JVrzkPpaXjJozRAcv+F/Kd/hIdEeeJZFpRKa8Kvt5z2k3cEeQiHcJX/R0B
Cbp62et+f8AOcgE/h1OvbZK5Ahh+scx56xpU2KhLnZVMUtFpO4B6TayAFytefdegIAmNCWlfsBqd
b2sHBnMgZlHvVLtoOS63zMgZnZGbQL2S745juoHvq4y4rk3+nPqhdFqZO9o0gtHa3gNGL4/hXLzR
7C/nbyu4kbO0tOY1h7oYFWIEMyVC3m1mL+pHQhpDaoU9KsWBBsAfUeXcvbrPQ1UlHvsgHuvJsZhx
HfPeNSUDO+tWZZqNS39ld+ukQ5DiowH1QoxDsYodh/OUBiSYeHwCx+q902SIXdPYw4GpL9QIADS3
G5CPt4YA9VwhC3R/V0IYr9T5sPril9aeVHvI/DNGmuW2SOjSJSSWa/8b2BbyP62Hn2qfeGtY2Wk5
vWiE6gBs3RZskpuozlFL0zwJ1kz36DAFDnzZFZUZflDJjN74Mwb3omIn2u2Dts/PvsoSTsaP9D7A
sEVgb4LBf2WQCpzDHAV7ce90qk1BXtal7KtXQeeEL41D2eJlAEL5pHkJwgTBwn30odZr6Zrrdiso
emAdyxV7IU5D2uQsQgrBhyftnu55OnsNgi7QAFaC+UA/q77hafxHf1jYgMfnX4Dgq1JrlCej0mjf
lkYKj+tUewQq8Cei5/CyXTZQmU+1Iq4coaZukyAjeYeZPG4seqJUAsrUID6cySojDtoJYZtnE7r1
AFv5xOhGL3IBVxtp4ultanP0jmQBnjHh5NeIpKnkKYrlIUldyZhw/jSIWWasAgq9ceR3/XFno7rE
MohKryhRL3y90crCGgzd97D7lJAU0PdZGIAfzqQvt/+BVZ/Z2JkKUoqJKajIociSFSBI19El/he2
KkuOZuaCK238C+lZc8R/FJecUa2k0FP4FLs4lDeVo2bHjUpo3Sq9dCp3G1zBA7xyJJ9AOZW1zPK4
tGtZJCemRdlQZjWfBZb9q+CA3NwDnX7I8q/agm4Lua20Q9IPw7uCrO+3O1XwwWWKB7DVLF73JBGF
YFvBpvJ3lJ/q217a7LJmIiOLnIET9sxTwOaRIorSQ1KqWo7MMLTzHexYQ95xMyhJpwudg+7e+Qpt
+/ZKz2XveCtu3jLbRQ3QpWX3eRmJKN+UurDavuKCuOKVktHZmq6N0zW7qyVWoUsOOLdDOT/zMdYS
6WseI7Yq59I47hqFMGxEneAhoxp5VcvE1eHjwkeErXD+JzTb1FfmryN8IIRDM4RVIU+vsEOjf2Oq
lxl6ohvxShxnLZApLERjqwnsdrqqONMejf/3oKudpNbnXVzFnCUvd34z2sr8hb/Y/naxdHALoYY9
ti3dtQjGXp+K7IvJyCwoho2GQodCA8EhLPpmOuZ1CIMGNuXPyNNe3rgdN4Lm5sSgWGB9EakKs23T
xv1+yk3hfiJ/qNDGOvgZkFaEaq6hpkT3iULHSwzaOX0zzmsbCAlcE+aHiL9r0BkcV3hD4c6FPpJq
H2WMETrlHQOYCTLyadOUlbLL0Xzz0G5hyGVc4WHj5h3sDhSJhuyw9Ifkjn+bVWMRFFK0LAQSvowa
E0qLk+3/zbJFs1QEjJK3R/5V8je3tHE0KogsaiVSkhZPH64Pa3qKetMBS2FYhKcyxbYbra3zWDSa
CcM4M7Gmxz8ML/zl73HI2vVyS/CAFROn4i4Pww5645wWcKDCWehYN+cdEoqPhifvsmLdgdtUwc0W
k4kmoWGzTZFGLlEuiBp7ShiGIip/KAaNOun1oiHc4yy9IKZagRjklV2HjIen1Qg31bE9u1aXHgKJ
PuXUgerYkUjVBsIW2z1Zt8JwMhXuE8Hkt3kiJrLQoBIw+xOoXxHuMUV5PCA3HZNHwFmOXIb9TdAe
zlxaZ3Uvcy5FQwwr63vtGoKwIuJs53wFC+0M4HPOkUjd1gg6jAGD3GJmOCfUW4aj+SsEAsFqgYsZ
uZHgXGIGgimOWGea9Tz2aF+opV82YQjbTSeqaIjexuiLHW9HlLDM1XsJQ9bRXH8CHzkMj5kybEGD
4sYKgYfjWMvB0zhw4YHyGyF3+MHw6JxHqZxS0ntQAb1wuxBTg5hidFhu3ZTy2W7mtylCa4cFWdTB
KxfBI68Y5rvZD2zQmG9Syakm190JEN2WbCP3RoZI/vRZEtqFxdSIL4sli8Te9BOe7/XMmHIW50af
tnUZC/fdf/+NPjV1C4r4RlI2EBcpBfBDhxIb8cVdI2nkJPpQW3RTxvyx3KNimJkMWOxoqnDQYEtk
fpi/qTDvXC9dqBoOInqus6qradOdqCQJSeoy/h8Y/+Qsg/xMLIgUeQzoJooyL63TPTz/m1as1yoA
LQipDyud/paj5CYEzWgfnsPK7/pJNKjwYpuutXjE2eI1lVvvwLQ8PQodzdtsF2/Yg6OPaeArkqdj
4uif0xH69H1OLJrvntQU8IGxkVmKaIfDAEeDs19C7Abdya33W23yJIf4EagsWIiFAdbnj7VgY4Sw
QBx4WrgGwJvew9ra0NCM/dT4eH/LVZo+bBLZwatYlsRMECcXxYnwBOJnhJbpMbpRNb11EM/IUo4V
hP7tuuUh/vzqtiT+hxvpLdXA31xTsXKS670963Y4gAkqQLsTmRqnTjEQ13uxD5+9ozvs9cFmYXv9
IOr/UVEt1ApnKWX5T2zRX+BORHLLNVmtlOj9xnI8LmqUdLbIrDF8ZHE8p1Ye9P5DTuhSQsbtrYsM
JLRmjaHGQJVA6IhEW5i1bgaPsyMCXRR5L6+B+ry0wLD2vp1BdyxAnjA6Q9zosGpWVz4qWPj+hfUC
wabJUBs7jIir0dNOIkcyIvBSPPsxt4CcwWflImmK5r16hikM7wzG8Dx8EHWyIkKDK/gfLcu+CxRk
1ugvkrf9EnCFrmiI9uei45ypKGnIAGd58WxBJciAgaA2vXRewQ+f1cvwISVLJOqWXcF4Pgrvm1b4
VETzLv8BgN6XOdfB9O871JgDzNOgQ9+qhgCc6vPUXOQD4x7gG9/LBonC6vqezSEMORdt+q4jHbP/
PFiiunmzL43UVx41l8+jPs4RXJSL3QWj03N3K7t1ASunvn1BLulefAUP5YLI1gUUchHsFvR9sBTt
BLx2N8t6W/yDJjtwBvArHXBjeVTCa0gwlpDW3ZblJX3gKUWEpDzICDljnWjQsQ78IS8hLzggFGnl
HNnD6ut+WTRC7EgOOhege4C35GjBosw2F+W+LWh8zX/1s8pTw4cjn5o3DgvtgRRZnZCdYDdzSkNU
ZZMryxzv98XxqpNyo5ff1gFhWt+8cK5pJntCFYZnv2Gaqd64fSQ44uD3PRKpF8cOniWvEdBIAEiJ
jPjM7fQi+ru555k7VRAArB9IsT8CM5/9BVkLrFxPJYI3vc2hO1d245bJHVB28A7ehk0UjpbfqCG4
+Md0004R1/rIti7thQdimZdnyyzwEozkzr8MGbcfOMquLJlA8EXsdgbE7RoP4nYpW8w1IIOlwyJ2
27KHmOendYyJgCycuFvTOZIjpl6quX/OWj3vcVDFp1zC6FmDK4emIUO1xLV9juzFYzyguddT9DGW
GbQ6813euvSAauqvBtTrUrhFQMKktpmp2sgvhoHT8KQGYMWdR9NWJ9vgW9rcahFrTS8OyMPuXXVU
04TfRyUZrRMAV/XUL1myCPZJfY/wnNMHX3DsGAQUDW1c9YPNBFg/u3oWesXXzmu9ehSrgQmZhcig
V2YaLs24awh96ppjoKVfS8CgRAUUjrPlEAaAxYqyVtsnJN/nMzACwCh4s3dCCXi0AW6zAqP0BAXQ
AkdR6DMF8q+m5PIOW8EVcOtAJlOxMX3WM/H9VLqzZBv8qEn7gUNT811sb6BcnxHh9MSlxVviTk00
Fp4PuWVirc7skyT63mFTNvj28HcrjEVF3cFYreGcUzkKdCntywWdEe7lPw58sMuH0cSMAVx+Kbga
ImRpE28sMCtmA5iz6R2xZAAKLl37qn+3AKAWJCxDmmYG+1QJbO5EQTbNPAGqr6knl1OKgpTjgQqD
l7XUF2IAywzJVAYvH9QGdtTG5wF4ERFIB5b0fLh3x0At9zc/sQmaEfjKajaSMqPpWHjIaMFpFrbE
nohhmsGIsS1LtdhwHq45yFMzS9ygFp7VfJUE93L00XShhL2yBrCUc3iPJKo1FF85KJm/b//Lx5fG
qzYOPkY5TJeIQHfMMmqJ+S0K8oAS9F+TDcVXTHPv0cQftink1mSd3LULXuMoAbTQ9rA6FTzcs34z
+p5fO4guzLud+BVkIfUvF+rq8IZRSfkhxIpd0AE+tjS3LN5mVvyUZNL4/2c+ADvkWWQIcPaPrFLD
LPSv1/SCbN21vv+W2MkGpgcq6el4rjZwarXtklAa+BgxsO4G+M47y1WO1PuSaUO9bdk9TQ5qyKJh
DlYZ5EkB2oqlepXR+9rpOEMZ1yFTsC9t0yGaTpu6SMrUtUVrw0khZzt5Zyg1HEJ0Fgy0yGb01r/G
t6wF1KZctQXdDmeZry+GKvnxBbRjuJU1NlW5tJjjXwTJ1mjqEH1eyd6bG3PwYd2XtMJTp8NaPSkd
L2NuVl5TRKtgWKfDh9ql6aiNu7foxF2wxOkZNuUIH8r1/0qzSffXr1cJN1x+RqKZhI29G8U4F/FY
ywCp/gNpU94Dy0gaM/6290BWZkE4VG939ENUajZ0cL2Ns/T15cCCBGomv751Qp9bM7CdRKEwGb3n
SRrED5gCWxFn6HfiCrTBq52o96uSFgPTWoviMuCHm2Ae4TIpQfmsp/h3BzzBy/hQtDuz3KFR0+mq
TKk944AAr77BhLYwugB4fAMT0v9zY2e6M5NiTiat5uDfW2HOV3HMys++iKl9VLQWAxB9/71BbnlP
CdBBXK+tBxLT7b0O+e7OILprP9mCyxnrrmI3u0SUTbTpxYgRLSKSRGU+sJ1+h+Jg2/XTZ+0ke28w
PKUMRREGg1/cDWovU8keocNwC0H7L8rsUi9gzqDEy/OndPwmP+DB2tfAPPZMCxVc2Y9PrMeZz/7c
ixz+6ilfxlCzOP4wyLPfickd2cr++ku+tX/rieLcX3xmMKy3XWvuv6vvpLRPpFkeFdVeE160v4mI
VkBAJ6+zkEYtsztmHiw+bKrwrI+wV3Om9W/CeQirbp2CM9w1ORoopI30UKi5v583hBp9OQV7/pN/
P8BEBlHHxpDt/SY248W+pI9Oko/R4SiamgTSUgFyUI2HwoqKapIpN2f3d/kanB6L8RONXD2FW4Ft
FZ9B898QkFgQZLTh1B/vHmpTeXPZ/AW52HwmCgLfeo7XrEIps7zZ3qx+vhjD2ll0tQsgGQNeNoer
H7rXY5qB0p1xmZ8Yd2LYSI4N4pJuF6HZpuZUGwXse+yFE+e67olxxPtawdsCM8MrkSYGfNMjPowy
1P5wWoV9JS/OdjQG7CpGho8mGWSrXxYGXv6w31pRFy4JHg1b83PZlowJ90zdWwY7ywlgofaEgS8/
+KDGPFeA3rVH0Isf+oYeS9C9Bl/24Q2LmwUY3Pwcd85xMYW1XQPxDna2XZl22pwPiDqvh9dkXC5n
5nGDmanAtbR0jxVV/62DXNKYT51E/i+yqfwMFQ3mHXg2Ct6bNGyngC3Z6eEYJ192LgXZGdxplCs9
CUt/XeH63SS1W2HZNJUcaACUPB0d+4JcvaxVxpxBJ9GxG1oXVg+lI8pc9kUnWE69e08iyWZzVtJE
vokAGvqk3ZuCybGlYRdqRpKfPmWHa7yvxKMAr2Fld230oYNf4nQBEUZ8uAHR9Ji23Io2EDba1iuZ
Epp8XjSNRLbEg5z/QenA0g6WzhU6LHix1iRMWtIQXTI4sE/JFNDrrqOMn4HxblL8gMGJGuaQE9bM
pQ4l8aelOg3oinjYO9PWNYY7aL5AeEMGjZjNdlfr0z4t/1Yj2DGhWaGNSmfBCE6Vteack+aQFhos
JapLh04AHHS1JZn3SquaGPoYc/aEH3qY2mR6QYJD1pyjR1CSG7wb+jh81/zOl1LyPj5ZmP+HzM3e
qbXd/m0GJIkb5zDqRzJJwue/CRerE10TKrYKiBNRDlV28NGS4U/T2JbAywRkPQDy/ZvHQ2MBnaNo
mUX8oOxv4OLM3jqa4xbU66HBU0RqzbpdHffvn2qOkxBJHbslV2GZ1pIVOYOEkAnrB+YCZ6EFebkq
sbPuu6R33EjTBGuKfNDZKbohZPl5TJCOWygS2HyHWtUIWamnAm4le5yD7SICRvqgb4aQ584MqbX1
djJq49G91NBMS3fUWDqf3vkEqYS5pb9TUGK4vhB7Vnl8FPCdeJ7skeNhC417z6dsqfiqS1yMCfI0
aSMXExzN8DBz2VtL/FI8BmTWr/LzY5JUgrm/fHuinHoCH2pdfBeZv7GLdgRWlD+gSMhmDcN2Jalp
iSBR6tDCR3Sb578B5vM0Ju3UAjp4zd9pE9sMC2HTEmfO0GZsdzmlX0SdNNFRvBfDlgaAcaiK22C2
Rge0uthSQyHy6y+4A73KzfG4Lc+h0zPwIH/vd0naX+FfpCIdB6/qDVkqPXkKkrs3bnxkEWuLrPAh
ZxpxXqsGSDh2bqIm41abscKRWSZGG6Uafm1Oip96wkByS4mnbnQU78AdfLLaV4bkTwgW5TXXDNOq
XGN+WUED6WQ6wLCygwJJpb/TpyTs8M+JMkDn89WxUgtsvm+ttfUNfLuxc7AQ74Z3Ze2xoPQNxu0R
NlZetOp47Na0jMczEJYXbo8RecnbRgsITG+Cldc7by52DnSQ/ya6qLCrWaxfZVmghYYzXgytveGe
r3UTAl7antLT5A4vamCJMn1Z7VRxaPcI9tYl7WvdanuavKHbnxm0WvGlXBCEbC28QKo8ClJGgKql
vzUDvB97ivuN3utsNehsO+nlUiq1Zg30ABiXaqJHF2YH7VwvH4u+fYO7dRzlP+lDWQLQeFTOiFfK
xL1Lsm73Nb4P8Iy2l+pkp+JKleZ9Oq2iX7koD8u/Zs8cYPrvXeiysS7MhobKp7gZYiZiYzsvlZup
/5dOer1EnBJX5JId/7/91HVGnr1DfbUIvKaSeaxhdvu32sRAyYIKy8onbgR+I5yq2oyUAjyHC3bH
/hlzX3/SC9c6m0vHcWc7DOdqEet6LN3hjka8rSEo8ObJn9mh1auLlo9gEOwACGn1WhKrdkA+7caV
iN8pK3/xyK32tcz4q4J9ildXzo3yKLYft6DXzfHD+ZYaRoM5kZlKWmPrrroTkAu02x9lbH3/XHHt
rSz0NqPEWcyR7Z1oKShGvHks1k7x7WdMU8Wv2aU0Drk6YYwuJvhAXDoZZdQnozYGy/cw5kXJtgXN
x4mN82Iq73VPvta0Uih1lpQGJKbkAfALbcdPf16FfwaSrzz/TO/8767c8LnITGaappt/eBciDVWf
1BZj2PTqys0ygBJR8IK34oYOwqZFXfQ7oPIejtS/RCfe4xIFNr3jjQWFiJpCV5nzsLNpQJ2kslCP
GOBk6O4go1DKWJhX76XckiCZTu2VJzXF4oiKUUgVTroTjHrTOAOAHknMsQ0rybwHr+V67SoD2LDP
BS3aA7Vzk6Zd9CPtJtbk965qdDYTcE14+j7TWDoNlrUnaM4o849I8m+mglzSXJe0htuGrLSh9pCh
rRZknfw/VnPcfN0r/K0OfHCsB72FEcSAgwGmUCSHJ52+SVMIem5xgziyfgJz9U0stlnsrtjSHp48
ZSOELhBr4rmbrPS2iLQVnQNIPWnjhCdBOJ1CKySCqlaUARNPK9BAot+EuYEzMcv+LGMo1HU/5x7n
SOyLZXQumTv12E+53wNifm6FwMAmVcHZQJDM09gXtrZOBhNCbpWctRzSvZTMjRYDY9uaGYRSXW+N
7qJ8RLH5jOrtuh6AiKrg3HIFhtnW1PXhEKLhwIr3RS91z2r9AzMgkUF4ve0pWKhoIT/Stjxd0BTx
Csll2A3o7t3ODK+BXN0N0bBwGhGaTLMsuJh+0EvUebDc/8bXcX/S7gQTFOHXS1vqouc2xRlpoAT8
zrOWR1LoNOj+Bk/dO0MJLyNspYMh7pQkb6v1sBQZTOf0tTBZMZySE4VYFMQABxmTUs6ILfVhpymK
5TP2iJ6j7ynt7QgzZ2SJricMy41MBr5KIXJyej8JXgiUOQDqsvhM2RkzCuHIc+fWhtbInCcG8pWD
mif0/OLdmSom0WnLLYjWBbeUKvH5n0BLvnjMYhYbh3Z3QflXXr+53ariciUkQW6ZNJWykjCp5ETx
7gx0CR2zn4QUU1F2hdaPyiZsm8ZTBxK+1ZUvIFJNd4CA25xgYoXIIq+6uFrDnhnSQmdeRNY2eqUk
Omzj85UgI6G/cB/h0tFfl5zFJPCAisRnFuQQ6D44Ln+wLvivpxP38pJBHrkzRZ0gfG/BSqeBD4O7
UPQnYshti4Ij7kN63fuO9TFESrSjPgyugRvcKJ+rfbT3q19+p1Hk3KHcoENd0w7oK81OSXQxTlGv
hyX34pJxOFrC3BTkmVnXL7vAau7iLUqJcHUxl+aWkyjwwx53Enm+a7/hPHdtK5Nuspwy8mgcZVhh
dQfaKtZUPu6/gxFV+pYRyS9JhNO5FkS/WT80CVoayjMcE2Ecd3EAVJMFphkKplTgKGMR/7NG9iq/
gFLhr4qRJYLME4wUt/0VflZf9LRsBcZ4WIdTsvFFN2G99My1M6Z1A+bObBDRz8WbpAn3jddPFvt+
1SIN+40+q4TqJSuTW6s5is/5ux9VyMSLFg8i9CV6nHPpFinCrcvE62ps5hLsQlnvS9dz2Q+Tq4tO
dU7rIn4gaLKPDaETK2cF4vSP8pD/GLVgLxJqtjY1QNaJHvnd/3mms69P/9i+Ndgna0o28To5nyYI
cSunO0uUQcQq0qVLd7tca3Ux+vOHowbBOiiwuyyQ0h42Fvafr2wp0Nwyx9cK3EpHGBVPxLA/S8bk
Z3cKlV1KgSjEUNa2//lI9eazpP3Wz1WgAMH1iw62nZ+dA1ZS3ut8fT9MrhYQ7ySg+Dlani3kv/2z
Ja78NIVLrYKdsFBp1Fwsn9Pe9wH1Jkek2/c1kO+195/22LU7nJfQmSQlUeaiCgQwYj3cVdE4w2Hi
JNgvyWOjQts8P3gCUgAKgJMjAF2wQ1ETU1sKsyJncxftBhN4g/LmP11rHWhARjUFW4hJAANzaG/f
vIX5q5NumFaHmHo3ffcNHQocB03u26nYecfEYEZIeIHpP3XoCWw+mm3YjnHoL6UYAoIF0iHXdPoV
ga6AZhUrSNOxpfxARC8PIS6HE8oEj4CA+oLMgF3s47Ep57xu4FRV2ywjSArpgYIykRZXgFEEGKL/
f9nIMW3R+Cto60JMNFgk6Q/NM0GXW1ClUZEe/ILy4Rf/1g9cYOE7RDqXpNfBmHQ/6MxUBGPVfkPR
OgLckc97eWbhUVxgByD1LfMVZGh48n18J8PCBrjUoA9WKQMv3lg3mGf4RGCsX3c1FNhwL1EPp05w
i3KOWefyGceQGxyI3njRlPGc8qykCuiVAgM0bFck7yhp7gnGXRfcEqXD4oHwXRlvFpMcFoR+sYcG
OSt36dk7XXMyLoeEaf2kPIhocg+iyEEd/vdaQPj8k2Sa57uxY8Xp3bSwwACJszM27miaT7Meqyci
JoNgYpD5A7pPWjga5YQr5zn6zyYn2YyU7ctqUlN3Z6f7sP71clLcWJcAMWeM4GLYmLJMPbLQ6OVK
Hjb1kUVAiOSq/o/O0zlmAMOgjHvb/jDa4GhBYlmairCiaILHrXkq/qN8DKhwUkl1HCutNbQuxHMD
0LrdvBCmxhx+Slxbu6tncdnzGw6a/xPz5itZWFz16+Utp7XlNChX10z/uslZri+C+INrzotmdomT
oWF0hwEHSzZ1qZuE1b+ZaphLFzBzE8Ruj2a4m2EdRnU+hR0npuFmCmsCH0FGILsRB9Xd/eBX67Hz
vHtN3mE3PO2rpXF2wp7K2ZPNGffNDcEJJMfbEJtr2c8Cd0xcUBEgA2thRHb+lyo+6w0PB63BS+Jv
uuwa3iSZniobc85hw7WDk1Cjp36pnkdRtfrEjvhn25hZjCrEH2Rl3iUznK6TEPUa0y2+1slUtID7
sdZH1meJMM3VEJcdRSYwMDpgzyRTtqpRFuWWXOT4gi6VdkCGznn1thihkBvi95BPj48J5Tlamq+O
6nikDDow1okPUf2zMo4+T1G7l28aPfuESG2I7jKSsIbxGRNw6dmHt7kfSpqaIg4M9PqunZ+vEkAp
HSExZc61H/wnA8b9Gd7gVnXeqBX7iej8LhFTpyyq/Fx8SjVYTK0dvM3VN7E5hv7Ow96DTFCmMEKq
rDwWcEAiRJ3HDLhbAFxDrCkPnsmo/JSrFusw4V/f3mqLSIHZOkmKnD5Na1BtB4+L1NUOi/jwAt0b
4OmUbUZtINbilCofZ5dGC5pzaXvwg2z1tgBnyUMHKUSCQ3h2IJLtqDLbe/rPjy1bS1JBAkeLQtPy
CW6wXYgNNYBSbms4aEnS4XR4xne4LIaN2Z7Au74EsRzvXl+7OP866p5JB9nxXyjOxbUk2xOpHoBY
0Md2Qf5OEH0QDbXeu3+RlZI2BCsCodEiUig23sT8Ky5MkHF/6V1TMlxlIZ8CQkA8yTUKcVpPiC+k
2BuB1simWFdXj/Ex4XqoZhUfrXZ3NWn8y8g++ui0g6rn6jtlP0EOnVEQpjBqoHQFJmhXCozfXoeT
NZjJUFbhuN/AZ81bLMCkphFTbX5UasxTY20VFF+NSmMxWGLFc5w2tj81R4zgPOrZWy2Q7AwEKQ59
XZsYa5lPpFNgfVCepUJ3PwRxxA9IMnyKSxMukfEpv68MKxBBaEvEUQIMKMqK40kAPNdUyt0goKU0
XGpyLzA4/6fL3KJs8Lb33htKUSz5ydCgL+Jgk7FHAnNanvND5cFFiAk6zoB1JOCUSQJE8BVRq44H
PAdKZ9cWc51UtCCl7l6PD9OL68bJ/JM9OJZjTf9y85/US1hrxbUFXU2lvpWpnAP+MmFiKxJwh4WK
Qwsvsc6pI2JKwi4h22BJuEiO+BSqTc90+lvP+RPnPQVRKDvwIaXEfW9Gy9wdGdj/8ZfWm8Ac3IzM
lGV0yeyE8LP8kn2Q8HfGxrBf7wXx2Ioecsmxv5rl5OQ+scpbM9V/ZwaOubqzv+c936xXifHpez3M
SDkPqLSpM0fC/j0dRzY8O+AQGZdMHBgAZz8OEy23Qkvy87xtLyUuRk94K1wC7JJyAJrkiiJYxF5i
Gh/X2TiHHwJaDBmGZXlGp8DGDL/cMS47w3gehmm2gjBxM5FtXWx6JGFFLuwOzwHTDLcBaXn0w97w
zulExS7hNjIziaVNvxW5O5SeWX8QTnjqQsYvr7o+JdeReSal2xStEAO4K5mQV4j2FYeS8U/GvaIE
Qb0nqXieYwqs5dpGJn+xrztzTg7EFn8d7PpxjG+0g2LxdmAY3TaYsNd4L/6P6tt/HeIv/XkZpQiP
/ME/jwGnYSrp/SG5gdh8TT8KNj7yjAyFXmOi1OqvQqsdXtjLhqsO9vEIV7Q053d6WzfUMS70y6aU
X50cVC7DEyRDyC9Tq8zZxc8CSUNv1UZXkp9jV3RBkJjMTlHud1E5lZ+DWi3AKYvdTDxxY0KKi3Cg
VpPc5FSFZ1sCBIcU4yPZ6XTlcoWk3kMxcA+ub4p2Kxh1LrVRXz8RB5WBkt7VnhZPVCU36oa4LlEj
/W0Qzj84X7T4F5gx5s0Zfr7drgmrWtNqShvagioDLg129LNoNX04Ciy8Oxwvg0CfWcDh1oqpd058
WunRWIdxngAmti7Tol+skCxzQrle2bO1lVzhbbwBaMidEDg7j8eR8xFr1s/SxGEZD0R0GDQUiYGU
8+V3RWvCksN3lxyqX+CzzpjP8UVFiNwvB++7ezPOif722rK2YCM6UcuFZJRH7GG+BRnsDW8eCCIr
FzNoNJqtORBNHw9lJmQgT993j+xMGEUwQmU1kmBJhrHSki8X9fCVJjg3Qp9GiYjUGWKRGd32iDxE
7kjr7Q+WqxAdccKtkd8fY5uUSMxPNnNa1bleO/c/NoO1QEOKL1KvQhCuVclhb8MEq5SamHitEd/P
/uIYRhEOmoVPYM2j19XCukVVmfVCmoYwJrwvtiAcdUiLEzcC/ouIaL+HVe3+DwsVACJhUu4Kx0JW
QHkvJ8WGhcAiupc/szOYCIBubuLhkfmXVcvaY4qYDdtqG4yJ+Pkenw1s9fGJPyPTUepTH28Eu2GF
TodqVpli/R0ySiuCMeivYJpfgYGtuPlJj13x05znzx8Uh3qaB52EqovCJlShl5xq4yApQTobz9rJ
EP6feyn364WoZB7GtVYJugk9281lBkXxJcE+du5WA92cuQRX6eawdR2I9b2kictgSoj3TAXUZ9CG
eVn3Q7lO9oWV1fJkCyJMq3RhasysdfyZjl29KVFI2xC48+I/6MAFUR+HGE45uV2IKpHmQ4T2sthL
6sLC3WyC2DtxZ8n8l2cbFBiJ6zGQxcstHl+5RB4U7EqFwdz/0Ig5S4L/JTftZ6CQL/L7MUHSNvT0
SZ3X/teDaiPAPMTCCF+CD/124+914XiU20qqWu/oLVRscvprAcukMGUC0ss6sLWKMKESwbJBZsQi
fiGvD32w4w0Und9k3eQUY1EFdj8UhTb69JhSWFGw7psWJ69p/7kqkzqH1BDq3xodsiRsWoM9LoEO
mwU8JToCR9VVy6Uok8ICVM8gcCuJVKt3KdzZC/a0AjdHu8/EAbY+f+lFMOgb27AYNq8HiTY8ipfy
vVvYJku9eQcYJ0WykxIzoiiArBvD2WWNovZ1wTtRxdOsTwszkXDtPPZMFsYgm283YkhaJ5Q9LaDn
fa0w9rqabQKYznBg38BSyw957Zs7knvA+kYk6ey3Va3JKRzcE+cf9Sx5n3Q8ijR3bGTZVeHT9FHH
qOELA4atzu/WVtJgN+fkyKUcQBOiiV4Ea+qRNz//AIMDjGT/OpmSZgMjFKxpKUvZ9fEqCSSfe+xo
93ZZ9osjcUSs5TdrCcZ7Rj4x4l5s0URph1oBGsL4ysmKZe2tc8YOeqys5KtX6YJYNKQ1C9pfNvEI
IiMQcS8JPpBk1jaFnDOOHgjATVHrTa7g3dDPm5wFYydu+XcuObm4dk8BBZiinWHf845PgUo75Jl2
PJhxEHUvXoSSEC3H/8z1OV8zikDA8TapTp5Efr7GErQ8u0I6VbcP+HFjtzgqFpLFtFxDSkBwlYTu
mffN2hDH3wF/c2Do/3yF5ZfRZDr8L024zeThibo9/L+WsJ0+AmpI/TbN1P0AU6jOhSECxmmn7vcO
mhLGk0d6S4kmYjZkJPOGAwIV43PQzNGg24SyTnzd93UWpJN0eMfPIuuNegKqCb8n26UZBNWh8JHM
BNaW3SXue6pk4xOVTkga/5wRSGHRUrC3RMPCBLm6kZInGU/2N5NVpg/StxncPEJDgcMXFExMqYdm
rB6TwsW5Bcqyt4iRp3ykwTG57IqgaiO6ND00j3b5aWR8ILevLR+uo8WH0w9LsVOzKZ3X4tklY6Q7
eu8XVmgvJbg1X8Cisu+fm/yInZEe1ofcrkDCnmLnajDW2Pbj2O2Xk6K6wzYC2ClN/sF/U/LiXFLT
ml7DtefJhuZqJYTxAfBK+k57aesM3pJ6tmeywr4HAtqiMCJFwHaRchMdyTAGvxcsTcn2DwrmEvnp
g2t7UAq/aRxNTXqQdohbSnbju2tOZwSnIxdDOjpNduRSUxguTypEVQ84YuVHiCpHdQqpl5pl7OOm
krp9VYbDfoo7Kkqc5Tfpl88WXD/QF3wdPnX8WFmqOnIHs1E66nW+RbqjmFYoeYUg1X3u/0bWn1LF
OUf0rohPFAnHyC2HocIoKLCv1LXFgp8FzaOE8F50qDh/rLN6mWXqBOIkCnufi55uMKScCDnH2KSm
mUd3aE0X8Y+SVD3eMTU805B4TyfWp5MDMPmnd+hH7mbnBObqdgqlcyrqhLwUNPPcOypB5WCrV4Ci
20ks6tC9ZPbaqqDTAssQtx9NBsWre56Uq2O8w7QtyOFNB0GSBPVqugecN6b9p8EBRRS0aCDfBU9L
uE6yzXtpPZjkNyJ8T7ltbkj6Xke1QP9nFmitGTvE79GQxi58kFdsd5MioK25bQcHzmpJKGghxIY4
tYOY0yfb4DgNB2INTMK6uEds6ZHuroXl5RdhS+YNksgcl0zOnLXHB948BAFk1nXJAHSHhhTdUk5F
HhPggcdC05TAMpnmSnK2Ehz4NAGH8BaU4g6XM2MbVCEKudzBSIJQJuiFlyMsb1qA2mftIL6nqzsS
P8fDWfLEECZH1VY/WeB0dDPLiaiusWeeK6kRgVMevQXaq42EVMLfFqfIBFzI0mKAYy9EE0ZC/naq
ilDwr3/P8uVTYbL3ITHBn/9lyrjPY+R10WXZjR6bZeZh4Qv8mlUZOwnn4BmvwPXjMFdxHEmzoO1b
KcF9hyIsTDm0C5Xlx8YLtHeUvGnLrIYmSclfi9ETXIg7ehjkTUFTJ6TIwhk4w4Z6Nl0WKnJOlDxe
XNe6ak1oxo7dtlsGZs2oV2AS/xyU1Q5BNRFRbhIxs1d0MTH8d82HOYQK1AVvZOzkvNF+b9WLwunb
2II1STkaOjwxn2Z9r8HF2nZgaJufd28M4mFzYAjS1+ElTwmjpCH8GaZxJJ9Zc4+RdaoX66hOCVIk
zJjfIg2BFg38IuO6hLOF44QEOFj6U5+MZXog4ydL9qn0a+Yo+Sq++lvp4eYb6Hzzy28IlY2so4Fj
5FKvC4nx0PIGuv1fILyIJ8GrBshcSfK686xbIZ2LbDP4Kea8kPW845Fqn8FV+H6O6uqdntcWhWIo
6t5qFtAi8rxiIR4mgM3FKvC1FqMSbN6jAJfZoVQHK4NjRGej+OpZ/wTn39pyLSXGRiLlcxnsfDm4
znIX93md2wGF90IKwDTEe4PQjgNpZkbGqBq0SklKNKs5//Hmtep9nGDhJpx7qtcI/OdfTVpzxFx3
MANOn/XiTzrGqqCCo7Zmqkq7wo/HBJze6yvS8Aew+ytRym1jxtWRIBWRLujJL4PZD0r+FJop5on9
kCdDwxyZl6F87JWPmegwh741iEMIIN6g3Vp6oqhOXAgU3P5292TaD6SBO0kzujWFCo9tVT7zPonY
sMvR3WmxJyIYNgPoI6f5EkS7y1CYL4rCnJSbB+gucKqT5dp3w4uKuP7BRUgEZ01rrd+5vqQJjiOM
HbC36zaUJ2p1mzBuxS2l4Oy/WTWMWzx/7jKVmCKZoFt56F+oh2i4Coo0bPVz7X39ApJcDPwn9vTw
2gRcpNKRlSt8wwzKFLwX8JsNQR0dm8hfmF3XUscn/JPGx5fzDaGf7/gvzyED4aNjIErRKVHpk+oP
xszoi5CBy2/5fQnV+1OtYJjzqGOJAhrckjPB0HlEAzVvnkDytE8sc1jmP9cRXNXeC77evH1l0y8h
8ESS3THc0W0BxbsThtzbuoS/wAArg2mp5PjzNozes206lL6Lk2oSNPNeSSKLaARk6b644OvuWQKQ
LkXx5iUZWrn6pko0a4SbrgtL0Aabh4B52tobaQk8mAogjVX4tUf5m7/hf2C/F/NG+tu0gK5DHIb7
pHwpebSyJIZUE8NhHZtUeqqXXXpePQZwkP1Ggn3l4IZqPX3d9XnlMXQk83TS8On0Jhfoz8VP1/Iq
SprNZGq8/LY4kA9mOLq71LS22pj9zFr3JyFoYIVkb8nytm0q7jHiwqPz3XLX4sYfjGo830irugJA
Su+nIdhxx84dV3GhqX+DKNeriWS8TT7Gbpu/Hy44d6U9TjTJuvRX7CMzPsUUnmzMRb1O0d5clJYe
x9fjfBqquyIJiOCm57tZqeSx5496j7qePMihtm95CPF3vtGv9/NhfattJRyclFGBz0iD6YViy9XB
p1X88i96tVFhUYSIrGFxZTQ9bqihxjKmWlaDlH8XGXv1VysPKC9W8kBkc4Q/xJmKvzhWjYSq3kLk
Ky5ge+F+lE7fPeLw1t0OgdZCwltrEhQaw1PqqFaVSaajpYgaYJLf5PXJgzT0TF9hFRSztltsQT56
f453E7Ev4j1Zl/RR8IhzxuSpU+hoMP7yknirSINh6a4jhuMxPSdWQ2yI5CVE2AslKaVz8dTr57oU
RzVG11bLe+qg7YNofYdohYRSmrlnkmPFR1jjhm8ZpjnpDPC2A8JEA0BhuAsLBvebLUssVZPY+yLL
of9AwSx4jdJyGL2Ek2cJMNTmmk8EiinVvAlWryYeKONCpJqGjSfXF8LgP1KIIlXw7pmvQFiwKfnH
F/5SezvIPD5S10NJ58giLBGN+Eo3ro8A7G7+S/Xyrq7Y7YhMwdghVT1gflEefm87LqnMZapelCGb
oONJxwFX4JcfhQBdksVzXssdYY7Coel1L/aFoFFm0WZuGc2DPcFF72KTqlLpMMqe44qQbpUpc3Pj
YIz2Ce8QM1+LWRPvOmTn+qi7J4/TTjA45eQd5Xy+k89HDb+wOoF1U3hU+/q2OvdwZc7Htx1g/1TP
PvDZJknIvOLxX97XFzNDO9dCdK9VE/JiU0bWxvd9Oxzb9nRr6aUyibHrdxWW4+XK+MR5/aqD4x4u
ijSVZrkgQBNF+DxDbBmRm1sQsz5eGQ94I55Fc/nv4QHBoXxf0qXY/sc3Bop/BwBoVkGT+BVt++Gx
qGw1ZLn8nOoZN7Iayrfzg1NcoUDRGVwZb6tpIWxew0ir7fH4gsx2BInPBa98i6078Fv97BB63AXa
nAfCoa923XqVSWrxbxdwzHbtz/fNf7oYKJf5Fw7yocdytxvZ4LGh0AZ6JD6UhD4IiLbcFYcJZiLR
wmQt8ZS0N0dj3TUGIo+RzqPLuwb1b7c7Hi4MEiKs3a/PRxn/yqNnNfrFMCW6x8sqvcdivYh56Ovg
fbSJ/gkgQbncn7QEjuDiY+Zq7xAW14Qy1Uvf8ds+8Jcmxne0Q3ZSXnVf3Ml4u2aQEmGmSx+XVCEl
S3X6sm+5UhEy3k6HzRR3OYD31+DwqAgf1i3XXISt+ktAbvC1ibrOxRWNp+zRzCv7GZrGlR8Swgac
vbMafd48PDp9avy11HtSyJC9Lj++BPDC8NhIoJGqou1kUKtRj63OQF87NRmE60a7jKzC38e/72Fv
58i06fmfzysu9La0WiIvVnUJNRsm446rc1Xu99sYHQpb7+z9AIXIgr7Np1nOF0B4UaICcsacFq9m
YS+KAKPuLqNyGWiW8WAhgs1SbEWRqE9NUQpJKs4xl4PEBqIr4KZiF1cWu7LmvXFX8Pf36PTBCRgu
7bhvYjEpAz5kSz8QYePDW23U7ZEdYBs/fLmXILg+JZsmG/9L3Zjy7x1KLkXxdEKxWiKa/LD+Cfg7
szN8e24HBKUx0nAFPHhMEMt/3TPljISy56HGMYPeDF6QO2FtgFx+Jri23XMUGQv5QNIXfGShAoYr
O5t2TvzIFzw5EYFopVgtK7u7Dch3lD05zfXIlxSRq8T2mfl/+Cr7xl9rpg4F76w19UDVkewxUxYZ
2WF6fa4iaHAMmNlJochNjtKsiT7bV/qeHhfNOBr4Tb9R+q7tB/68tJc/ygOjnLaTQo1F5Aobaf8x
BHG2U/WYinWqlasoIUuut38gJH5oPfskn8rvPSqFRbeAT80fsAdt742eDBHlkwI9V+Fy3O6c0QDA
1e4E588RKbOJ9VQ3s0M8Wcd1FQZn8Uox9+IkS0W+f/L9DQ4aRbmVC0llkJx+XKJb7aZgxBor3BXv
WyoAAXzj8/cd1IdlyNqF6gwwfEnBoph8wHZW5zBfntIU1LPCvH6VUC7Z0v5ehHyVCPvmZLdDyGfO
CaO9FVubBSmBMh9KijhUOGT/tqxv/BvZdJvXpELBhLdWUPq/pb2df5rUSnv3ZIuLtOjzOP7wDp2g
yAAeK72uRiDFVTvQnXHq7qscyDnU+Jl4Tx2DZvkTBY6/p3AIWjg5P2xKeCu4ecVhEILMe8zbP51k
tMrb4/OeQXZ/o+UHEZ9MUKWFZE9QrAgLmeAEw2XcvopE0f5m6ZW4LMMOx58BiPV0XLMhani1D/hJ
6GO3Tmhyb9kj0Z47wMwxUnEcQHA6ui3BHdOPDreurApte3u7SpJpmzuElsUwLP21/3N/9Xpith+o
42IzYxkefk3kJcEVeHm1Vc25TGu+5+gUXHq2Nflawcv37SHbUxqDjaTq/1/HMJpvHhvGUMsUI8/5
8qIobPmj1tOTdPXQe9TZNa88rRD0IWrmRW6aKkValEy+QB8OZUhQVN2tEZLYFxreEGe/jXtJRFcl
UirvkWuggNec52cfUDkt3s4XfcKWdco2ipd5awhkjfWbIIcvhbF/DG+HJoH88cl0ydDbaq5KMqYh
T5lIP7jHcI6NpoKQGnoutJm5hSeh8eGRHkPdLr11x0TeZgDpStjVN0rEhQlhkXxK8s0LYaE/HJg6
7aM8FQ4tsQ1LpXyWzFZQtHQ10SE0AoM6CaYEF1+b7GuGP3gNj4W8tAwaJgauSRNR4+wrXgQ/JCn3
jLSu6BYEFpHlCmzuokFVIhv78hT9Q+MS7hdFbKyIdrLjbtGDsIW9YUnOryOXlfsdfiw/NJPwgBDF
fnHuls8EFXLmiPlht4gzc3OVmx2+nwmowPMRArIXjjtJwrEHdIBXyQp8u9qZLEpVbGlpTi0ddiyt
Aa11MXD89j4iBvsxMIBDVSjZ4y7rFwOw6CBGmfHvNMW32iezY3w/N2AKgrKjLkAPoxYMH6j3OzX4
Yb/al3FlUYy4XJuYsu5j355ERAaTIP3r90R0RXCXO9ZZ40aA9tDu8uf7GmepoVLm+ktKa7w/568T
m2tDJ+ntBeH3I00SMW/PZaZ01ADFC7vwuon99rtnYWr2p+oJAYm5TgoFjUYxRQtO7/KwivaMOp/j
zQU6/q1zTYMkNdbeRJ7QdwRK1RkrKWBnnwpWPEXDomV6aRTOeNknED1O/lHYW/m0p6A3dTHKh0XS
nvUDljPWc5EyJ0Ylebn7UShdEyl8I8FgLwdk4ijNB0XMJ0Yj+D2upNs0Pi0kyHLRPSDE2xclcaNU
VQj8u1YWtxWKye5h7x2g5kYrhosvQXuQXG3JCho6uw2U+Ld0D8BQapB7GL4uBSU56rM4nD3esW2v
hmGVNaghA23+EFP/lz2maPrIEYZIR7lvbH0zR2wrHogopma1oLaBiatKgwYl5w9aD9JnN1yrmBKh
KE9zHgI9N+3kMyfmzIdKJ8+h+04xskkVSFh8wfKpAR8dijCADWG9hVQuaKel5pCmhbP2Vl2M597O
uTbu92134qp2h7apCx0SqybDF4XeLl8PNjpFqyhM5SmsrYbS86+c0iC07J7pBBqGntzLCGVZ76jk
oi3HNx7BRk52pmzfaH/l/wWg7dPH438WkJgnKLPKK2KQ8XEurltUGUKIgoQJogNpOcT4fndmGakp
iGYg6sxFt6uEIKh7SAgVM4L+LV0f8u/CMWy3+s9qB9c57VU1JK/MyNW5pEAy4yvd6lgh/BeE6LW0
zN5r9z1b2DceleqK6vM1g18Y+L6R+1jTjfTVLPRzobCLnAZ8dTa+VwhXuJUwzOz3CczZUgE/B7qH
zvmAiXzF8UVLrFI+TGj7OgPGrhFF9z2nJOElRqLihh19i1OIp11ajS6DJZYGX39PHQJOH2Nu0hvN
9D5RmlqgE+T0LcjvJBLl6eftxFipLxytiRahZ66Jmv3xzEB7Vpice3VjmERVnPOF2hU7plVRnAzr
CkMhNCRQmV0vaxsR5FXM1fjTX1fRH46z1c8y1UUKglkpQxxPcPgh1GBUFPnWav6gPPiAF452YtDa
spe/V/akf4G1H3J5yo2kqXtWapjiv87+9UVVU7B+OW16Q/K4aU4U4EVPw2gd+RmMC2l/MdubGyJ/
duvVDD7/s4JWapNDlG7AM3hCQMlMvBKU25BBrNXCnsyEBllsQl7nlisbRE8sLBiV7n3M08V7YNHt
AKgljAicAgB46rPnjqhYiKVZPXnMmYkIfXljMn/bonSaWhpbXyOn2kG7nvtFKAZ8Dx1I0KDKUVaQ
yCsEEs6kJivrZLvoNALyYksBebeEF6xG4JtXfE8PVbXrpF92+2Oki79CEQR95wjrKj57HEJuy3E3
wzgt/vo98btE8qG8hVdvRfuUczql38i1oXmqUsfQ7eJf2PN3h4MieqQxebqt7eTQkfBm/tWqy97z
n6HUa6wF4/RWpQe1shAXw2afBkwV0TqRcCYr0GQO3ElofghNsRhhQPVKlm7M7gSvKgwsFhQmGwXU
A4YHxIdlBrHG+qxvOlY6kAt+0aLROpYxzlH1DxRzLNW8Opjz5zf6/ONmLJ3W7+kvy9ii7E97LAp7
5ETOwIw5TFewp464cwhFC3mlb6x0sI6JLjROpXFFw0F2R1idO4TC8nPaJucULlJWEpevqN6E7y+N
zwdDksEo9u8gGh3bqCwYy3asg/DlGa0QTImL/FJnyKHuWrPl9iLths429DhpZoyMTY23mW6KJgjL
oiUmFNmqSRjU92DGUg4uLL7H8S7f1YprDUIBBRb4kxHamAHf2GsuWsDnw21BI0NJ9kbqqcuBt6nH
r+JPlerr2LCajjgihFfGH9eWl+cinudODUSjGQlswoildBkk0f0MOAgzrarjSZGIzCdoWpvskzK5
uOCMLBSawbvzgf6UxLQrTVe5wZd4kL0EnNlhUFLgI9T4IHm405314C5gGBrug72bwtBEclM0s4QJ
FYSVvEVm8sd5Vsy9buVPt1PPQQ5JSOGswE0BD/Hj715bRNrXljB7Z6EmpD7zlNPqVFvXYoxoGYQu
ZdpukkXyqWAU5CKtUdo/oZQWlA4W1gGzOVl/mih0HkdDLpK+X7mtNsGe1RI6bpxegU3+ZZk1FIG6
qlteLfAVHBkjehxksSgplidZ0VN3SgjgIUTaZwvhLp7ukVjF88/LKjabBk3yYzUqAGOEGbP/Ztdi
8s3unV88YRgkw+bhTlQ4gedk59zsG2IiZe2pwzjD4TYF+xrP11fz9YpjsTCS+OowCI9yE5afERxs
swwrG2JzHxUPyCsAhQA4IV1FW3b9ot/ka2thg4yDhtwHJTQkpp7Sdf5fytylqp2gPeYCao0iGLSS
XNn7mr3Gp4EXF0XCwjvLE7M+hG1FYfxLgE1zZ+YicBvIonExIj3oAD/QZaPDG2y9BxOkhc7W1ODh
D8PjUVC+XvA676hg8YxBXqTxYlQsCJ5RxP6LSNkdgcdFdH0DVLRkNThpEmdlb0lo3hY3EKbBybAd
YVUQESVcv1zw735v2zf5YM6IiExwe4GCiZuxTbyiWHLvqpubmvqRsJ67d0gg6Nz5iadUQizXuAe3
j9jKn2g/eDyEkPLf9KOFAIepSPAH/mI89t3HZ7vE7OeY5eQOq58w035pdPvlacSRzTlM4d7zOGq0
sD95JPbQjgWgxMTChRl75F+o5zaPlvm8ds/YvoPWpUpaiLktomsbsW3DAAxiT+QO/Sv/Qac88DjM
8K3JXmUVS12PyP0JFFs7+WfBs+NIxiS//+XdSsHjvoR2S4AFkZI57c9Fc1YVr3zmMdLR5gAM2gtq
LuN3mdHJNf3lH59n3c3wtaQx847KPXtw5o8BnwXNmMAv/afsph5NEtYQ6AMeZFxsF11l1HScfnbC
1DkVA9+nwJA6wt5+4Eol3OMk2KVQyhh5pUdlecebwfhAb2+1KR3+9WA/TOeWqH33zzSrWcNul/oH
ZFG6INdX/K0Fxf2QzEf/rolrku48NYcdc1RiX1rVTVXU4jT9jtPwOHKLw71Em+Fhjq0DCDxUjMFB
ZRpenol2Gq4MVHLh+0vlUbkfNMmZfJUg1QCHz8RigPMp0PGVQH2BEWM/7P3DMiwUkWJ1A2DwlXMc
psWYkQpPY5UoBT3QmDTane+f1EAUG+xrRvpmfs85FhpgE1LV/PNqVpcoL3J2MKxiePQPYhC8RhgK
FE2z1JHRj4p8mZDRh3Xnl12UjkQaAO76Gqy3/5ZjduEXwh2EH4aqwklaFb6mEDmY2BU8tiRyzbyF
TFGLl/Mi+woZLN77pdWr10LaJq8Rxceu0eWkmBWV+1574p5CtTYbn2TtF7yJRdrqah13B0aTggFb
6/lf6+zZuAbUqJKRTzj1y6mJ55GY8KCzT6bIreYJTOI4Aq1E7ctWv74k6nmRtJN/ZA5E4FPjgrUO
DQwrq6eFKUqJSK+AT1shAkD2eDzyOZlv25R7qViNNmYaDYNKzHDsasDZfRXnGIvAS+qGM9Vd4TmP
NQ72jCg46sZ6e0FaRVE4Jbj4zQ6+p9uI7SmgcGeo9RXGUxDkwfuTZYOo44qYmQc6sgDKbnpYcvNW
VttlSIzg7xeHIu+vqdQfGWaszsjRjmLpxHGxYX8eYitZ03ELJQZM4UN8ix9p+NzBneaEJLse91jM
29AWe4ebhBN7sbiDOuQpppjqXBa+F/m9z/g0WIJmSoEA/CtwtCSNeVb3hMyP2+FhR23wLMq65viR
YRsmyoJBa7UWgeRULplMhirSZuV+o9PNNY/1tTLnY1TxtbuDU1Gj/saLNpZk3NErymMkVAIp6a6c
Ew0spT2zNdmbIsCjb03xRnY4cl7bg2XQoYMWT4UkY9rXxWxWQGIo81yKrZD4WRn081GCK2Xa0TR7
SJjK7WTDYfGij46E79YtKqvGBGd7UgQ3vSw3dkWat24E9II2j1y2uc6kSS9ffiV4yAjIPcLOATtM
iPHky9p0ZJBdiZwjmBCjjinlUgUWksZ0JFhnbqkzDMhs50sUl/ESRU58tnwL56YbiDBG/OuKEfG4
DROagmH9F/UMYHF+DMPKCC14IrtOtt2BHbAYnpoKEne61GNvUVQgyN86XoTlFvntGmXAJ8EYkR0z
GM8YjHHIy38b6Y8cwBmjajHtimya7i7PKoqHl53c2u8ig2geGl09Uj9efZaCh+JEithivbqdvATT
dZ/dD1LQiVRESfRoHUtdY6w/fyjhiLZqLZ+7XQItWs0Qse6iSnpOGocqzIMeyajIy+G8zgWq6bZO
w58whVrjdGylUKFRbsAe/MeaDgwYNpgYEzGNKqp5y6XRqOL87lrC22xhXVQVcEX9S0qt+COTQLJj
TY3oK2Vem42mts0AVyu9Fp3WqAzaq/V7lyHoD8Kp8OUEZtIU3R9EHXF8gdIdeQeSBvRzifZyTqhD
8NHeyCUSNs24Jo7ZElD4bO3UCwLT4arjntqTUMhmFEx7iw23f6HLsIjr6aBeyNuMQqYsRlhGovFi
LqRtZuRVOB9vb4rfPZtweLJjYKeKoRm+LQg69ovi9LDTfYmOGJGFHe98CkjgYAJlu36p4Bpp08bt
HEvLSGzCpm4yPcY5YlED9tIP1TqCin5x8BIwIeyHXoAPCNl64fmp91vXADwfcr2yMzQMJHHQs9K7
41z7Xo9Tc5Y8Y4GQDVLJIeFqNVWP4kDNdedde66hqvj/qlSuUs3jtx3XZN3K2n8YGYjqBSo90+B1
/kM6VGojqUbK/ZDsLtsLlIPCxpysbf77f57bTJ2ltuuh5vwcl6POrYKRAlj8ij6SUd8s2QyVLJhI
VkJgLuqd/tXprbLAm8fVvIEamWDEICT3UP7zeUjzTwAKyt0CkzkNG3tJtUrI6lviPDghVPs6fjlo
fNIZ/LISxQkQPhcqmuK1K3Xo8XzWqAWjvGG4Qy1kJs1JJp8qivzWhQzxaCSLdK7jXjwC2ZVweNc3
2O45t0AQNPzVxLw0fi694W/5AtcSzwtdGc/JjIqDrb1ydufo0l0CGe4botZILGF1QFw5ydK6N3rz
A5BGT427g0JJvDuZLHyXmWwcBshyFBz/jZ/zfmdIHZejHlb9VXU0aXhkzlKdnjmKuefGR01ikPET
XRCBuETGkGr68QW/IbCcsijRUN+QKeBPCqL+lFR85CffmgsCZvi/INOZW0KDcxlZjX/NP6NxrlD/
ANafczUZzlmDxr8XC6VybRL+UxvGy7LzgfRvEu+toB0bO+axHaAxgESnjxLLoeqsWwUQ+AiI7qYK
B71Q/WFlE+N3dctT5q91oZQgL+uYfz41IqT1LAt8NksmtJvcbV3kZfnEyxMO7ezaVffArMlLWUrd
9UDE7+46YmpCIMjm8HgwT/vfdVaY9k3FtTS6tv6mcgHkGZZMylrQpPJzi6GXtvbAoqi96QEY5mjd
EJ/cqH7LLcaxtmk4ATMYxE7F3E9XKVETpLaJDAPvRn2o7XB774lSvIvrGfsluIgQ3pLUhVXpcBGJ
bv1jFpjO6QaVebx03nayCKi2pctdPUTUTH9UsAF7u/9r6x/FAcjSKRsrjC2MzkygTpO4TT1Fl3gY
NYQ3+eOMr0CE5Aqj3QBIHhCp2x07iEuaxZIlZZkkF8+Qzb192s/J3Kcq4D9jL/k3LAiKnBDfEXLW
mtsSnH39xb8OH58Pif2IpEj62BUawc9NQvyy/FYGgtPNxkCVl0dVOrjfbxynvPwpgrrueGS3ugiD
Eye2w/Zz15ijubIPrbtB6XagjwhI1wU1tniYKYSegyNO1i3yE5NdTfkBEDCba8pNQ3eBt6Ouo5M7
Taz0kkNejvkO+gwLU/HL3Vj/MwtwrMwvAZsY7j6LM3PW5bzOxXaHURlfuxVJN3SOZhvbvsXbDpk/
6oaMqpUHxY1oPWHLaxygp3YkgG1Czmmv/j3a7SYgyaJtoXUJ9B2Acwc5u2RceG/7fi8B6fWW9+Ij
Bu419QQtrsnQhOiEXKsqg6d4nbjijpialE/LFnzUKSBj5jWP9MrlKiXiIX+3VwtSwLLK4sRzlSQ3
gSYVXR4mLJQmagVJoYrqFMT7/ucUTqHtd9qDysQ/1VhzSa1K2h+emEEUiwD+qWmc5K7esa2owGKS
oHn9rUpsf3kBgUji1oYANv+puOWl8AwczgV/znXhSwkvZ/+Mj/4uLtZUCj7c7F7Ea4cuNcp3laBv
FKeaN4dXjEfu97suZOnDVBdIHsAj0CBnjowwmAm7I7V3Ga/Hz9I7EssN/v4qhahTC/HCDs9V5NCo
ZaUUP5IzwXiT+2ufRXk9CmC95FWAHq857fQQiEqUBd2HGbrGqz7u2A/DJEoykRkyKl3n1BMmzP5e
3hy7LbfxgPJ7CfYY3puygDvywUKekvZ2shb064ee7xw6pr5ooeY0qG15A4FxXkmvnOcaZsZzi8Ef
x/q0ZAFJc8aS0GCOl/+Mz5h/CH4TLRn3uoipobcdg+CtfatJL3B3gzBVaaJioDvBExELkqQ2YUI4
fQsbFD7LDXpS7n8F34hnbfA7t7pbpkJM24m2S89w3R6FxQSdYjhsmXAA+JDPFytqN/y+hSkgTCDe
gJBHhz3RGIdmHsQ0e194rB3agN/HaY+Rcl7u2aicOdH9K3zOCGYk0vJlLHCSkYTpFljgmWsOEznF
zRvKmmSLp1xlxyCJ/1qoB9Fibo9q2KRXmdMxP6SbYGG/0DE5wzyYCCN7CmRCUGGdDq5i/43NNGgK
rFDXXqx+QBWz2ynzmr/80ZDYOb6h/FMKYEB/pZaOUEVD0wfulMoAg3ATVxSW+vO4/bqmZZGTHKAw
q54ZsMELtCv98K51iOW7Ev/6+6a5Uypbc9tPan7WMQkBY7aebN7vyIRfd2aVaKtYH3ldvWUHwHgv
Pp3etDVdhIewvzbOmJmOAQMmYttYLt4fpQ+dREfrkws94hPJlR0WgZjc50MrWnx3ceT8J4wAgiAa
fX9A090kwm0LQwP3qZlsFUmgUM3VrdU30asVoxcseNCYe548sBAZfyWZ4w+2mUnIGl09lGBHRfI9
QDdhVeGeVcZ3hVvR2/P4UYOms+kg8uF3nW8vSU+u5MIAEEhz1ry0DNv/cKt4ReHXGggg+EzsEhb0
KEW+jinPO5a5qwwQrf77XXg5xxEOchOa8Frf4jzmiEcDkV37vcLHyR2kszJi/r0AuQR1ag+T+HRQ
kspY5NQJ5Mj5kft4OHzC7K7OGAVw20kr8EuWo6eM9y0AjXsA8fr5pHOuUuwvTra7jEhheHrqrAgi
vA5/8ofapUstvIBPEjixYrtB32GL4/YGV441R9x8GmLSHWO8UMSjM46/jIBIzqcAP3mTzBw9vG98
78x7CbxZq9y8EM1tDA3r/S/9JW5AKjTUr0ST3Y6ArvlRxUeJN9UOWr0PHFnMr0afiXYRa+tpOnaj
9HMPQh+LotXRt99zT96X1Cdb9MUiZd0ASqg1bXiGiMecM49WngwUIzodq6/zImwRtJagirgt5VXb
yIIlkg9PIr7sGQFvEzYyj+x6l/+mWCcKe3tOEftWSg3yDNF8gtcobTxJesH0epxThb/RTaZKT3gL
oweUJBx2AtiRR3yXJ6bFAhQ0gBuKYKfL3mf0e+qhedUXebq8yZjA7/Ex1y092Tcb2h3D3GWcrMZq
wb2U5Gse5ad5AnUzv9NmyznMskBut9F4TgK87Co8MADnLXEOExtBg8NXUYoEudrHMdtNoSGjXmzS
8T7PbVleygXz7WrsaMxInU08I1T6NlrOiqZymCd5PD+h/8gcsea2FYV6UFjMAzY4Hs4K6uo4+FFl
LyKzulRG8eI/wLfKxPLPy/SJniqpDltEwhElPdvHrkDCxDIsAOmexKjPQ6+MVjG17o2HcCNMOPyw
3wGX3DqXLOpMQRWZBHmJefGn/JNZj3o7bkHhLyFv/SlXA4lx/zQv23oXgnB0gz5AHbNp+mVlZn4E
1F1dUJ/DiyFXb7Tcx8D1gg1HsOWFdszqQVqtK67Nf/Q/38HWP1uJ/uOGRPAxDLtkCMJPQVbz8sSg
2s1uJgUfPGL5PSOmBL5su9mxqKCEjJVzzkl6bgjI/BYsj5CldBRHoH7dcVALVFGuQSusm9ECtdqb
6I2I5CpBfWNvJ1yPKClZ/z8UVYN9dOUAY9JsDnSY9QQyHZi3rpXI+3TJDYSeMO0/L2R4j3Swwosg
YYWHtZu03yf/EV756VEdyiVtOtfTMQ64ZJQhKJAbrVE3iU7AxL2qRuwxkSSWCZLb5uidasSg/6Oc
EDVIEOOnOuCrPVxV6ajDGAj+tAy+PKcsqChY7gN5jTaMri8nlW+4reI9YCQLAybCO6vuQJwkCpxC
BWzwb+W9DSEMzMT6UAg54yC9PCGuZvra22V9T3LFmbj9JDRcyqWK5vEEZRolMKNP+5tRAYVo/A6w
2KhHCvyNVjajENZuCu1WvVwqnFy5et8DIQyhGjxJphjX0G5ozKMaZHTq4r0Wsb0J3czbi0I0C2ns
eIBhKGO/KF7ntT/cdr4P47jcKrpwW1wZ6u5H8wF1XS7fQVyCmdzN4XYlX3VLe6NuCkAB9uaVyWze
YIEES3h6rYwtp+V694yqtYZeaW6TYC67I23QQeI2DIGgU1R5AV6pYwx00gHi3f9dava/cpQLsENJ
g14momSEudOP9ReH/vT8nU/JdS/UHpw1XIeQK9BFk3369paNxnrro+d0y5p7/KsdxdDxavWYmpQx
usNe6A4IEwtKRVsH+jxtAYQV9RP5pFrMB8BevD53gkayhARKX3jbT5QaqWnl/K4qOjd4Qswx4GWN
p6vy59TYLiHtBfLLqPvZSGw30V34L5rqa/wyCthFDZQBJDOEhIXScmSNffU/dYnmCJQmjAPjSXIr
kQwD1pqCwKSxZUb7rCq6ilxz2rsrmfVtwwsSvp7wWl2EOZpcAWXCNEwshZJNYT4UiXFtzH0KzBd2
//PUb8SfaysfGvo2D7LdG5nDFpOUxlKZlW32Cs8rg5iMfkuFffq3FLYbgDti8CFXHfRIR3yfWzBZ
YX8TEF2VW/iVu1n7EzPbWGOBjvIMPuUyxDx689fpyVfq10O+/dfPg7TkEaoxFwgSBZNy3h0rAml/
rTc+zPIr4HKkTvYzbSu5+yWa4/Re7I7IdrYEzxyxyCTd7ebV9TtvnyvrpoVaoxnyabWRjWvCga8O
57zVoEMo6Y2MCXicjCxQvu/MqMXu5iQlf2Rhxd6w0LeEVrEBp5Gd1Hph7thOPkg4H7W45H9jI5Zo
Nl9akbOrJix4dPFy+DY243EkItx5Mf9n34i8LmpxuoJi19sf6uMQYRnXB4gkei/+hi97n/wnVC/L
YemSD20lkGzBbD/AzvCTr7NDWUzdlD4KSIm52XbYzRzFiR+qZxg6c5IXAeMwIMSzp9ud3Q4fmQak
YjooDLUMWhw2i1KCnWMmg2alES2NBpgc3A8/WrolQTJKAYiLVFsUE6+sXjlRV2LH9lHLC99lmIui
kO8Bv4QOM+92JX6P//NzzU9pJBkJjswqyMjUPzae0Zo76rXoTLDkJN9Xq4fn+R1WSR+UCy33quOs
gBq85b8Xj462wm8cgxAS6Q+AnA8j24WUivdQxa0epuzW0abA/MCU/7mL2rNK/oHbWvLh5KWBhtnM
AD2q/UnzSbFbNRTEI/gJEP4Wqx/tzYY05Iig2gh312IPiun+Oa8L8mnClw5oosGzMGwBznC8lQeR
+qb43jCFu/IebmBq0BzFau63uSBDTZTObiwWZfBsWkNx71mCQCcY5NVmyqq1KpszgYINvpvJHEsE
LaSu2Q3lxQEj0d+d2+OVhiqjH4HLSc5LSTXT4qqGNtO0OLV+n9S2Yf9qU1Lb8Pd5txUaakPf4CFh
O9vW/6ZyT4un3buC6o+UfaAIV9bYoTdZoiV9aWcp7SfMWnPpS1+smS/2ZQpJHDpS/kAY1ZOkrFj0
ZWXLJ2jOIs6Fha/q4WlnCM38V1aIwXjeCnmweHX3rItExIzYjpEIRrzu1vGRRBdaTibJ7DpuVSVc
pK19fWpxpE2LITpONcFFHWRzTarRZ6AOsjFgotRj8vzHJUGA/+/fa5GxWFdO0tKycWmuK0P2iH7G
xVVvPfEqyZIIyxPOEtmVuVCDN46Khw4MSI2w1I1rbI3w/BogcKK1yCIc7cGa/o0Ie/bt2mq4Q5bN
Bks6Dx6pbMRBYAiLplMMj5677TtrGfl/wE3H/xsx8EFOiPL1suYYUud0TNUN/iak6lWmqjQBKZQQ
83BcDmffjbdw6ALpyOZCODQKhvNVtHxepljuyRobYjZJZgVxulO01Z8B1LKv2pih2gxg9mBuy6km
/FdMKxATrgikSg7qvctDz60a2Yfcqpv9o482725BXMAx/P0zuV46HjxqPF7oXykZ4/zaoQLGcSe/
PQcwrXeIeqhLQR2KC2QIcTtBQYeHrCiNQaaK5CLWFMvZJ3ReBvBcjryIPXvtusK3vtLHQUoymlPI
i7YcxWLpZGsf9KTaJDQ9J5Te5sw1UsBq+MhmrjhFQZqkT5uatahviZ+NPk1hI6zRWUTdePNVWGJD
mNaIJVlKc8vd2WqwycDTDbFPRSpYRsaJIl6v/3oifY5zXhromNNJxw8BuikKbigVgBeO4lyaizan
leoEZlVJwI/zZBAOGxUQChDMGzmhkfW5fnARVQIx4Vi4AgvoqRP8iiMCBN1rWSgJAPDjL/1bCzBu
y/6tHVwb27zXgRqD8gtDZpekpcdH2Jy+0GQ7Qo37RpiFa6YPBQO46hCF7xXu2J6N58+AyhQFIRu0
o/sW2XCA4B4OUBHNRr3wXPgT2azWemIH3yZyn6PIvTk+9d7Xq14JrINgYWnva+p2iOFU5o5HpD7T
nkKZ97sRmm+fDjdWEMDax543d7q1sT1Xg5pTVSnzchhdzUs2JX+/X1XSyjUUlCOs0JENsd0m8P5A
Uzp76k/KeYIcxcA712Kq2IvMcX8JbTwqH7EZLU1E+6GuI8zUsFq1dNHd3F++j1NYu157t7KZyHUx
49lcIkuspPIAt2DoUuLU2tzNglBECp6R3I5RotvoW7tUaIXyvK0MFbh6Rw9N5HNqCTGhg9Ep54IM
E+Itf4TovM1ElPeLZ60f0Qy4ChJmXso0lMzVFZ084FpG/yGD/vlzkfep6Umq+03ES3T3zcpHfXTl
DULqYXJB+oPllI1K4qVVI4mdjP3SYBUPZp0dpcIPbXls13pUmIEFmtTSj6uiJo8Cj6B9b/wfUBnO
xilslkk143FNiMJhFgWiHOlSUSb7A5o5nP37sIQya9eH4/nQx92QPqFqylwbitCg2sCH/FqrM81N
mZG6HaM15yG9QUvSvKAV+U3O02+YVe9nLR6T6BmFU0jgQhpMvCa75zv/bRoliq6Kr0JPrLsyoRzK
VdgXkAWQENLypX4l/lhSM+u+4udRyw7gpijoPRtYlD2SwRhPFXwxwIRYRJwX7mAMOJc/dQXr5Bx5
J65YPNZEDQT5JJsUtt7HG5q5WUtWKwAkzLpp8ZrxkYqF0pCh2fzgHbpr3/QXgsqHnpCCeiTMd+2K
+0uNP//5sgvCAy85KPHaxDJOLOvRYQO1EdeOl5a4v61qUuutanPm4/vv8WUFgiRltj5+sI60sRwz
EOY5YZ1F49iezxEqr5Xh7cRqDv37dvQ97Agyt/9tiiEz/6RnpRczUFkXritIVrtWWXGLegz/duhf
MW4c6PnDDNDKoz0nrS+j+P+GNmInAZuTaGoK0oXvK2arudjMxhW5oA0uDOTyvnit9gHML0dogMR5
4aatgxLhuSDRKANB96wMTckSE5xb0WEpiNBuU0d3xPjiUJxXFG3o/tvtGNVdmGTcBUMDMnENNKCr
O1uOeAXP1HT9JyupE8evEyUE6rGiPp257SIZq5A50fq5ISUeYiOZ5PAvqxxA00YgVNSxQTYFsQW1
kVIHJQDGv680dIhdTclv+LV/QSB1K/S92UUJoPU5WIvu1awKQDe7swso6AtkO1f1vdRT4vb2oqSj
Yda9EUyZj/mMclk64zPlg7pL95lYBT3tmA0PpugCXCxLtCuKS011uMiwzlEkTJ/90pd8MzBiGg1F
uXq6ubn+pU3aoBYnA84jhH0XNDhMxZXlTYxP/Y1fikiftTNM2KOPd1WfyI/NxKkcKI3vM7BdvAEr
wjefO9+pD2ThdJQaCbsvsZVjt3cFR8wgvFCW87YpKNqFI4AEkiDSTsga62XWbUOzpgl4iANP0o+y
CbNylYvQ6dRlkY9D0SC5vhMjVDxtFMV8Fzz+bLhRWUA3wblW0s0OfhZ67EEitdTeTdZeD6udw5Sw
DPivHYrE6XkP+7TfSCKp1uQgs1HnFvcEaVxOUKORXxVQu6ccnGfwcFVrf4wO6bWNFR9dVgaSsp0g
hf6ltdBuqKpS5kxw3MrTJiSfsmrcCVveoR6AqqBUIMzupd3VmgBTZy3JEWX/f/ggbvFM65H8vHTI
qtitCmbc9PiMxOEI1kxz+zTNWpV7al5SQrVZ5xamyKnkcz6vmpWS2L8o8+Lgbih4LbeW492vgQ37
wktZeXILu86ONZR8vlM/DGJSkQcF1v5c0NLGookT037AZnLAY9leGh6IxhrY37eYrqCTo3Sd1KWJ
kuvID9xIqbncMiNvExDLWPoUJhlZ6gbV3DZcumz2sFY+eAUYEB1RWRkAgtOHl9Mi+e7hm4vkXp22
Q+/M3CSsvuc2xDBsDvxqKCUqbGEXtu/x4TuBTWoUfBJ3mG/ggC4EuxoFbFbS0t/vGaELTxNbgFBI
dGLQoObT70lAfRNZDtLS/5aLjiudaD1PH/yZBXDv/RM4Xj8mbv6CNpithGo9viCWcZRZFrtW90vV
VC4p9GowJPLEKJLLL5x/qKf+5E3Y/npM6C2LWR8q4udj0pPj8Mcs2wFj6RCCix5m5lH9aLbaHcw9
B4xqIV3VBS/d4dX/BQaFzkmiXLZplM84qBAOID3lNjfFRgzKhO4ti+y/PKl44IBMuAr943dIhFHo
ppeulwxiVhtetfG9+WLyeIpOZP8KSbtQk/YziMaj+N87I8D4pi4eGmMJZWo06W2Zs9aUdhKjP/Aa
Rh2VwlULo0BsYPD1CXI31IJRaBkOdu1pS5c6nOzPPVuLhL6Hia8/izvgKs4Eo1c5VzY1t0dE6Yst
5UygJDwi/TY7a8YsHVKmxH493fP1HbxTiBLH+nacVcRU02ZVsUNaM36ftHagJHp6HH6u92nxUz2j
Zdqb1J/6LWFwOSVxHGkO2RR86kEkEXlL4YCaj2j7AkD0QxpwkGYi6/X1IoFc6ZqWGR6nzP31GjU6
yQU6IYlthwVSWXtUV3xrXtyqWv7DHuZWm5c4dIAa0T7mhBzKugMOopX2WYvRazOCcAXN1WIYTTG+
K2f+jn1g404Dc2LqiZE1jGA1v0oxuwSE4X6WiVzxWugN55cin8+aYGUkF2BIOLrugjLcYHw7PN6b
1rRGMVkPbpSasExvqUEMwVcKaJbcZM6BAYIkFCLQY/iXkq1YJevcLSXDMYkchAdJPK4Df9ToFyxb
TBose/mRDoBBzdjd7O7mouMipU7aY5xgYb1V0ZXT4dvYUo4BQZLA0sYUhrFaNKY7GzfKj78LcN2Z
cwSPDmzUFnoDaJsvheSvydRYycfKqvsJ7etYPSiF0heUJ7mTJ+B6EcAx7RgqTkG6Qd/cggBYrIqL
FJwME4P1nLQpWPqc42gcqnW0gopPuwfFi3+IrCWP3XB9Zn/zFpfneD1NbypfzDYmZDgLnNk1Lab0
fCT1Jh74ZJEGTmLZn1ptU2z3hq/0psXLZHVLDd/p9Axr5bOZzUjjGMvh5YGmX3bsq7f0pbA5L2Cl
vAUh8z/cYv34e71k8QjvwM+XWdn3ZE/s8awn5xWcnLioFkCKcW32lg1n88WQ/qSMQY4d90P/PQKd
GbYtoeKzBy43RlqgSteKadRevkFSkaLximJwqEL24iXi97MJaEg2iLs9QLvivCoChALzbUrFGMNJ
i/tKBYK/74mPSyeYYsMq61r1HTDKZkLtequ/OaEJEzgetzxh0hrtECxpFQ6ojI++sP+OHZBQ4+5z
lpEnDgKiR/L9Y3M4GqR5Rq/cZcfpKOeHSzR2XnvsvFTyVGG+qvM1Pz61IfC4SS6ZsPCgPAVFoaQc
4wKJ/yQjrmEfnyWuiPSdXfAmqHZIcXyvwJQOeAOWhnqvatygbKw+HhKq+BnyjiWQdPxqAICOVXkm
8rrgPfyt2595u+DhZcZrk991DkcXI1zV6UUfubIX0TCj915KbCLGSPF9AfiHX5c5ERlvI0rbmogt
oHpI3Fppi4iWjDkGqCI1JYT+k1uxMoRdju4GeRCnXviw9QrIQHzSxbqpYsqlBotnL9Q6IM4wN8/b
Vc377HVK36uC8mXVmdQ/ooeubOGegfOCIfsu3V2tpPZ6w72HYmFXGqvLnOLJ0MqvLpxyhzicB1Ra
KlSsLYInXfMUrllESuL499dMAWfzlqXlcPXsXOhVSc4qVpWfb5qULmNWD5aXR4uj9rCGbX6DH1D5
nha3UL2ECdL5MQqxNYtT6OuSNt1zW3IJL3YcfcoB1SyfMNbHs3Cm9TSqCDOMhcGkKWKc2VWrRSFq
moWfxyfrAdhTEVE9f9goZSb1X2qBoOJjrxffxzptBip6q9TFT1T7VFZe8dzuMT1qiSGVGOyqZu1U
YDpUQSRf0yimu8Fg4e+4kJbetsbMaXo5aentdMS9bEivj0xJCqQ67wInRrhwCDeiJo7HgUQskOjU
TrlaNZsaHGNH15ONScgEO96RdZ6tkjbKn2fUpZqfX4zSmLxo9M5aOsQHIgBnYUGur+63qJm5cbyx
ixt6eRKLzf3ISH3tx2hcwCWnSPy+MHbLFJ505FESH4wDCUmlRKN/Z03NMy4UEUVkoCqE5TZbskow
8FGhdK5PXGA60o+CXt2p6RRcHaCMFTnEE8iqf0MCI9buzmAEOGqDLnvInminy9KvlWxLJhlcHwIG
8l+4OA6Q6UMbi2oJQHawC7qAf3KYW1xGgg2uU7cQCjBU2KzfxFULvgeuo4e74B05OXo6AEw3erQ7
c1W1ZAg3NNBdkQB/J3Gm22H0XnE9+vIc53mvIvGz0QYUeAzyF1Ja+q/8pn2iCWaLE0TfOmVimDWJ
0TrB44fA3m7cPliLNerTFA9im/4yiIASNYUb60H5ST6MEQLGRYB61Xxeubo06WyAWnaBCt4BG3uP
7PTCUUeB7NhTfvGAwbwc7qX4Qs9ryqunVCShO62v2hv+Z/ngZ3ckZG0o7WJCfKCgkHjhwZg7sja1
tKSPiRxilHGL8GgfxEaHcUkAste3PCcJeQRwNOVDY1NQ3X3ljsdFs/aS99xtkAhn0Jpp5m8+RBFW
Gwnz6dpJ6dANSu+SAK96T9PU17lkM4NW7FuYHNMj68O03fezePK89kK1kVJy0JHqOUraQGcmt4zL
LuZ5T/82JGfU/EN6+uaK+R31mHHlX+U2vRpcYTlZs9bTZEgFk+r2nxZgj0vhJ7eBrnmZFdye52Eo
ALakSLCwlR0Zn3C40u3pdcbXr/9KosDNsIPnnzYZzyftqCZcVW+qo8X+IXjbgOVrYPo6puyVLj7A
4VkpaGyIADm6iM9THvpzroMJboXoYX+Vkd4cVSJ9l+AKOn4X1UDwG9gH9fIRsd/AmFODhPFCTzS8
Tm4/9nDvt/86WO9+FD1mVKbdMRmmdqBcbOEU5SaNmoJGYQXdt0nlgF3M/VWtRJSYleB+LLlOr0u+
bt5NCshSDblZ7pvKtbVvi7HoW4w3+aYTa8UV6LaLHvaYzHxI8H/+wi7hBDw3s+q9kmRp4/oSPWf7
9BFAXTQ6N9gdYbaaa0u7mNdbsskpZxH5JqGZ8i3UfRKR3gP7lvIQgzxlmtT+Dz/fDwuX9+o6rkzw
ixCzpbEpKax71cliYspCdbsssrPs+KYHr/GeFIni5wZyQklEChfqqHA+Q3DoFP+N6mfIZL5XT3e8
uMZEVqbIB/X6dsifqGalACO2Ws5VM5E1PB37cyafqhmLRUMkWTP3yTEf9gIJ3GPejKLX6ARJQAwq
4rGmpMAIkqfLieEW+uifYzhYsL7xFa0FANybSg2gSCEu77HgtBYBd2GNkaYLviemsy+pn3a62fJz
DzMHI4LAsZ9wHoK8wCQYBm6s5vC2KaL0rWEl0a8SFMd5x9S5+5pkz/Bmt5lnUYm1NTu2ab9KPBcG
tDrRJDkvi+yKPJw0vIZ5ETNtAuqd21zuhQLlxjpPcxKv4glA2VdKM1222tYLPEPTm03PAmFZ4X1V
WfoKpEINTmKhfeqUd9PhSyZErvIjMjoatBabggO5jTWGiplxWqHWLfMgQsQlwNqRCyaefkFfye/8
QHMdZ62Sijo/TBqbPebL8oF+sinmM7XQAsvZ5EgOD3O5obp4Z9ocZ08DJqUhbDQyCvrMJXPcExzQ
Mwpbzc2bcc6wcW1yNVeigdTBmehKhOCi6qsEAJWPA+dFV0TjK0CXvcwbPjBLujp2cpFgr+fawIb1
9Bandf5kRgHU5y0Mn/KdjQPyIFX3u7nnoinsnlQ5+GvS2C57YFExut3sgtabuoDjDproWUmdJODl
tOMzp6seW9t+jUPj0vgJaX2/Syua7qEgxnnpn6mhkTo0WizS2AF4xzdGd7KsiFR2aQX9y841Q7RG
XCQCibfU1OhJx5TE10VsPtTEtqMQDeka6GRNZiCk1lY362KHzfGMqRpJUr9MWoESYuE9S9ZpEEog
8kHO9I7DC+JMaoMn5UrhiYB4Gpn5S9jncJJefy6jG5BEYrNHoAHcwy9YAiUCFu8kQ2Ixlc8104tI
LDePbxNmJ2GcvRCjMjipuVdxaq2Br4CtTEtd7vfjVnwvznmEHMHre9rzsfVpxXIDT+l8Yor6FWK7
Oa/3fFwvOo6PVg+xfqo6ebVfkqoBxg0bYI3fjSX05qNeAoZjEBp2pPIH15bFKqVkvsGk4KKrAAkq
NWC6WnJuO+GXFucgF0qo34m0fREa9uST51+8+oZAKpdi6xEeRJHtFS3m5Vbx7rVC82oMKnbnBm/f
atzkSzjEUZIgMU4d9j3xPmk/0vFh0dJptbR4i7nDMHxrTi7D6HaJ4FuHYpsR9FjhVn6fw/gL4tLo
Eup1aJY9MZh+WVDh5PO7+x2PvQ1c17vblHtuDfH8YoOKJYnQgivt4t/m2E7T+skRo5Cnc3ISNk72
k4VJRjdUbmf5RHXsBwqkavyDNiwxLMitkGfuRg1GHlePUFGZLh4SG8ap3H9gZuudR/NwbUrUuKqf
P+hl32C9sb+4c+6Uet0ucadZ3sR1oVpnnG0yT9xO6pgogGnwJDu5jse5OipPy6OVcfutkJUEVF4y
qjlCGCGfAoz+jCwYj5mdsHi8EdKtgWwEd9fan0f44f/bqMlOWfEoV0iSh9KVb8UobkR6L4O8KzxS
Wzcob2EUyXoaaXLiFIpR6xNSGynxAsZYZJsPzRNsamfzY5aY9xAFCfCODhXNA3cTX4vw/ie6J/+f
AQGo323kRbgBlFetH7ev4esSahSIa2xwAYU7svajvSSjp5d/CZQRx9xinCu0ok7meoqzZpfdHVzr
vkc8AlSzRR9cMIZPM7eJ53BlUuQvMdqVk54iEIpISKhDWZgpQuq49lMUmsKGrCQ2l6JK+iLwKNzm
xKXQvrep+TuJsQ5qjTznhbbuedXqiZzObF6qSnBSUtJpui9ITT0C9Dtmrauhobdk2FVlclUnTHS9
7dv21efo115jBsoQuwYBWVNCiZ6KQwF/OTEFgBynzPnRMGCRq0P8Fg/mm+RkkXt5AGMqGf7qA5cJ
ZQFX2Zz5CqEzlTyyQFx3oSlH1XBl/uxcsZ6IvagLFHqvDLtFIPBvmOtVVi1xIrfqUxjPeca9iQVV
YU0VpRkrRBTYfL7RAhAjSQQlXERcxz586OdbRTzznChpGf+FdisftvAL4GlrkINFIULAUcqBjaYc
6/32/vrv7EoyWewJ3Pb6Hit5iLj23l+F2uLHL2Ifq5ZM6Rg2BZNp5ImWD8ON+GVEfiXkRk8R2AEa
2J+NGe5jpvdUSLjugZNuBGdNjE3M6gWedtgYoik0vBEXlT16BVSeC9ZXsMbw7vq429+99GQxDaHl
c/Hl8iA0R5/jbF5CtSAjZOiq+HQNZfUKpuNSwjK12PzMu/UVVBxdkXjNtsL1fVsi5S/5V5I/qQIU
dFZOpCO2BGeEppy6BS5oqWjI3P2nDNQan/Yuz4us18Z8EarJCufEhsVPTNN1S0XyTyl2FeSV26/c
8ozF1uQZvy1UWYTQFNVCtwjJMCbYiZFyEAg9p686fjkMBTqguLc0Bnfm5EkIuGelR7dD3ZSusuzv
lGal4CtzpHIPmpNHK6771Zz67X321nOP41mFPcjInXxM3XXCZH9Go/0pF0cr6N3RdDE43P4RtcsM
V4dQ+XMxfZjpVrbCK0SPnKI/b8F8QA2DoBkYiHwcYqKbBRXFiokNA3PqlK/0ZYFlqbJNqfGbonp5
iRMacawHCjvYt7+UU3GZbX11i1joXGz17SJLY/lAjaGEgf8ZUVNdBZjrHSf5dfyS9om9DTgFX/cW
HuX0uv9dUcehDXqehKfvk163xsgMCgZQkQM9/HjLBjxDIhUPnwFRVBIMewYG5zLjmdfflz49SEsU
LTes8fCPy5Ozs38OK0TiMaGZogUrOMGpYqFkoKaVMfLRRNcxdfDffxT4Og3bxqByTOVy0uEBkLyg
6wgekhtnrdfjWsp4I8oR86Sj1YkgzWttJpBbvcHnkZzo7Rl0bPB3v9TwRq7+VA5yydqC5WpddF79
bmUJnpkd3EZl3uyXcHKEzCplpJ45/lGqjGuTfpgzxfgT9a2+KhyZMf1q6ZQTLKFfl5Lax6Oxpbzv
q0Zh+DEbVqO7l3/HjjZuCglnxiHM4RlcCNHF9NozxL7VMBQJJXWXDWhAN9PLxD+uVVFEFm7tylAp
K/vnmNQZyhMxjwR6V0/Upa436x+iORp1PltmlI33zzCj21iR06Pv/VvbHBFnZNLl+DTlkUOlRXlr
ztNW0ifZP0WQWfit692AOXdQs/GP5+fCR9RRhrk1NFUK4pExWs/ZjTB2Ddl24KcQfXZxBh8Xp7n/
qg7jNKEYFEXIbM4RNbWqCUxMr1uhqEgSnFMJWNqy1tI8gEbvDvGqSBeLIMMti0U7JqfWiFNvyuRU
cYz9otjSho7eLXn0i3KZizYa6Sxt2ZhTVIACmZ9DayHB5NiauDpm3XW71mwlqWi4XFKqtu3XSFEJ
trxdqW3R6xEIpBrfrcyMv+R+uK54uPCuxp1Fg5uWrTFt5uvUYxPrXgtKkLbPaCPNUT1lNWKqfjlI
bprAsDk5xO8Z4hsj9BAQTRjkbUkgf1U7co6Ce8X0kJoXKuXIWHr25B8pNGWO6IVVDdcIr7668UVY
ZVtX5IfNeCqwpk23oJi5ucTDaGACdEbDXonLKtcsteIjwkwiXTyl6cWBr/B2GJg3UsfrksOF5rza
duBKzkIfg2GLJbNwLasiRDjPS3XBn3fu/5cVYVG3W70JTmviMFjomfEqCmPNBqMDqllZU+fiMZkx
Gc+MtlOJs/3PCYQ0BHqL8ySYaA0ycoI8QO4fuzKg31ywJQjHKfdiiMwFmBZ19sevFICw8MdzLGG7
+4alkG3RGGOnN0FnQGxZROP/BxCdfBHL++Rhusq5VmwK8kZSoF548/QE1Hr7VdQUF184bpzGyLSN
dF1n7FC/svr/FFFH3mlxXIGywy/V8qluWsrnK7Z84p6zkLIu3vNoJg5v2EaZ4ClnCyKGxeYx36gO
NugNB3yjpHsI4o/iBbT8mvIBGW+yI5HBlckOHNn0OJyMjMX3BiQlaalumHnDFWvrRgczgdod+sKR
3r9MftcoGo7nB3P+i3WWjklo4t86gio6k9In0sVOMgrwnqkHlKwFz1MmJanw0i566FzvH/T3C8hu
tNQuLKnAMjNugAzwFnPYEH/P7w8uDiv16K5NaGRRuKZwzXmc8H64n/j+jxwy1AoUn43u9HCtzsBO
xiD6p9fiIBRGKbCHhk/FMGlwvt1jeW01U2RafpSughpvSTZ3PcDICCEqIGe3q7Go+nY6CXuGXIJj
T08CImSoW4NOfgaEiRaTIGFFC+Ww+GNvdzh7KrWh81qnBgTAbvfI+VuOE6eGA8wyl6V9mwV5/6MK
ACTXX439CsVlfaw+76weoJQMaLd35zMsFw5fEWA7x1shhWbJZua7YixHI8bM1DdE4h/9u6LV9LNU
Eih+VF+kCMfpOaP9uPWwY2NAnRQO+qXrg2Wh1FfhY96bhdPhM0ChlN+Q1Ku+ETKlekBxpob78ODj
fr7G3P411ctZr6/ZRDDiQXH9YSFaOAdBnwLqSZsvvFr1tCTwzM8CvsnnAzI6+U1hHfZ6CeGDjPC4
1Qj/6jnxv4Hqa0HY96wA01h0Ll2puV2bHYRUzFXHS0aBvaU8PWP+4+aeL8Poe7lbUnuw8nx0LMfd
KSujKkWbTcLO50wrXgBViiy482x0kXte7MVTve7jtp6vTm7gk5WNj8VdS6C/FzkCST6yqI2lI8YH
fng5witfnOF6HdtGPwahhMuzNqcB6eHqo2yj3Mot7N3kNcX3Y5Xr0VW8g0L9ZnrnaGnjfDmQkc1w
ErDz3cQ9c5ok8bfYsPDLZ+Ge6yLNPx944GytjAIAyr6Gh/OkI/LUBMeM+wnRBvZDvNpH41dkWYCd
kWoQB1heuOJJDt/CUDiEaUXbgBF4PqEb/wwiOy83t/9YCiWwrUKqy96ocJtgHSOQd5f4skAk+4bE
azEeNU3PPUGZfnFlUGiIH3ZoF6Y+Y13H1oQlZMoBaEGf/xXGHukr5ZPANiPQ5LnKx5PhvZRilj+H
SzefndEV++XA/M9aaVUaJrqAuf6cNmw5wVcXWOSu49WA3okOS4f/7cf8YhdH9Zula0gMecg/KsZI
gFE/bG7rc9p6u3CmEA4JC0wS3P9eL5BL8a/9z48pvYxnewMQWoNgdyzHRrcrO3qk4f0NPqdHU28d
yGftkpUnfUCWhxBm7L2u8MH+nn02TQ3jRVrcoCgigs5v+j4SaIxfxvjvw15Z62drlOWjWLEo4FMr
9c8j1GbpxZV38ohwff8yGLjHgQcixva11ptqEjXQuN03sxGXVbJxFAsZMX8aUF4DX6sanvmxo4zd
mpo6im80lMywGI3B5qqu0h7v+SQijrLjbqTjfQ3vhrdAyR9eid8v8NqOLrZlZC33A1af+p/lJZBj
6qUt5WLuZ7n2zY77tiP6Zo+clUaczc0Je9U2ec91T7iFw4ZmbG9OY8JHZjF9xFp6QO65LsPk2E2P
VWX2auBF4bn7UcvB1+VwEg6iXsCIWlHbPENrjRDjcgq2sD721OTahhbnBdKiotId+L0jQkmBziYf
lyb9KzPflpqNh5SZrTwH0LoLFPUPtF7mgYIqWKG87b8vUG3mJuwksQ6blg4ZyCUWEiDEeiT7EAun
pt1D/l1dWYW+WIzoW6A3pexQth9yyXW87MTCqYxgr6q/kXvym/kGwXMKz97sP5joxWNUtdBU1/uZ
ye8+zAWOtw3jw/r46haF/bfEjQerNUsRQjxeYLTYhhs9gLVW3ZkZTygbTBi8ZLukMsdaQHZLGWx3
QympXz7lG0MV+13QGiw8GCj34VRbByrCNl6KHNioDHTa83lymSCNBsg+fBuke4djoInCg7pFRPdi
ocvFIE8OP//8t8V8wQNQHSAmq13AMQdcjSdv52Q4IJ+RYezd9Pe9d0osv6pbiKJqBjhveI3pDfh8
pjqNW1ZKly4PPBYFgU4ohEjAVpC8iooRqJzNrHvdFxK2oIG2tVOirq1NrwfpIIbylTLpdqnKGzLD
xm6tUz12rmgIB3y9/OIhZrSNF+UUd1syuQq1CR0CLM32kDi4Q6jweArRmt1uh8KkZhRptH2+1ak/
cDZ8UQCcndtehuud2txDi/QDCGP9uh12XmDUBMEbRKh41gnE+du0j0dt2seC90es+Qgxb3rp+OB5
1mul5pyP2Xy9fFBxxCp8PccPuaKfG5V/jvEPNCDytsqFRqXr32+jtO84rYMdoQkf1ZA1ek4eK7SU
8MK1+rnQISQZYbbOJPE8qmrHKj2TBKLKSIFulgZeSMNelmKzXEvep9RKTO5JocpIBDuaAqpLNF4o
1nOz2lgIHfN+oPfpAQYXH+iHTj1om/xHon9ohubulJJj5fM46OWFJFQncmif+hgpKhh52FxRmUIT
NzTnJt39GnUfKaI/GHF3mg99b7M4BpFRk3f9EBUrg92EwXPotNf2Bq7thgmTa1v4MNZVsqseeBqR
aisyGqB5wDGF/EaDjfb4t9v73L9HszzwdjidWKFBNpNNE14BZ5w8ry+b1CwGpGdRCzLVgjlSPJHI
kWnBSRL7P19uouMbMh7LKNzZhzHUDCKx7ZgIQZgz52U2zZ06pskfv/4i9gOy8Fh792ewrfvff6XA
XjEMaKLEcLjKVLPLXrwIkeEdKyQGVRimCfhxOC4bu+GEbrzK8mQ+pC0oaY4XgzbZVqPcpVz4fPmT
W4gWzzTZeT6r9JXe/WCMFRBG07uHG2xWmCFAGuY9EvhLy9yjK+OJCNGxLt3cCBoWfCg+0qBNGpZM
qCzatoNxGr+KRV3l3urnAcFdQ3TSQLClxovWREdmRsZB+c3qNPbDMN3mDqVzq3tMOxMH1xlqpxkz
bVkXZdXcjkUhs7zg5Y0006BVcy8EckkmeTxx3xriaYzFITwaEHCAKbadY1MesmTuXvR2jR3EUBiN
fJGR1SKESMczi0MYZXD3Bgf7eDWoley3wdIKM47JXpPRLklKHe4gMfVKehMUJINEYs8B94No9C/Z
9krFQHx0XyK66e5oM6MRzeHC4v/M/5HhhfpWstsSOwa+TULf8koF2V8yHs9KM/OjdqApmnWfjEb+
DSTvwZdPXpdO5xu2I0PhwfwMf9JP5GzIl6JtMMOGMeL0nTLMSnMZ58cQ/q3bycSlv5v5Z+btZ7vK
KD30D4Iu08QOhcc8aFmT/VqwrMWF9jtYFnZpnQ3nF//jwc9px2ZcrdQLxUmNGgkfDzQbdHRSlzVA
s7s7OADJbkzlTCqn9r+8VArYkSjrKU895U3fZMY1ii0un5IsqxWkOVf0zWxjTOEc6wRuUxaYu8tL
+YxQ22u9+IJRQalBirCKhY6ElL1aMjTqRXSZr6ZrcpHpNOMnDMjblRsoml09gZ8hqCEzIrqwMo24
yxKIZsA95ZVpUhwkYRikV/C1LwS0IjEdGRv/qItT2iRcqMuiIYcA8R8nlwMC7s3biJjfsK7Lkmi6
VfC7DY0ghL422K5DWAvPtKOgRwE9HSl5XWZcUia+Zroz473MWNhb3EM48kubKv7zW/2gvrdf3YOp
yYN6SYqjdGQyesX3cx+HL+rLaNbv4r0AjyjPfwO5zWOiohjUU8irejPWUiin4ythNerOvLCyWk97
wmU1iu9n2EmvWfdbuyBUURDobEbYSkyemC+gwMkUigqnlR5xEnurR+/BMirPswcQCMBPFMG6z6A/
b743VQhp++jZ0UdAlz0HiG7HMJlkR0+bZqG5cAg/0sqmJ9XNVqAqTWoSLf6mkJOmpICNzQbHmAQK
zgbKWczdxhUW/9fL1OoXISWreZXJEdYXVSMqTWeD60sF01lweb0DutfFwPoBNsE4Dv9yu+6PCpPR
ojRMzExEof1J2EJWQyBB4Ycu/kFukhkD57Y9oCCMz6ew1gw040DE+tIuSnMtJ9gD1ubxWGlqMF/j
XQu7vIu/xtIeQM6WudBcmfe8cAlug4zxs4JshKVLOqVKP5sDmhk9iGmZQgbPt8naAJhbnTlJkAYG
RDjSyKfkFKdk4sOyplyAH1tYfT4M1OKRqvVZLg4u+FQ8/EOc+H9GhMk63NmTIUO+SAtpx7dl3vxP
/Z2EO1nSylLCwsWVqdC2XK2ysq0KrsqISrRL5Lwd8JsTUZbgEmuZn0dj8Bm0p0iU73lupqUw3A1M
rZoN+xddILoodhSBbsOF53Oh4iYOQroWQzCuIsfDiUGCb2sLDM50Zs8VdcuF/Z4Dfrh4LdC/3Ozr
xWTNlVGxxIyMbpePQUvNWLFoT7wNBH9KULe79fxfN7qIiTNQv77jkUqYEEM9yabIogI6YP3/zZTV
KGG3RL+wtZ7NuWgF12AD/fOikrAcMtwyvBflkayue4O+94np/24bjjyg1zpn5jUjQiSpM+cUkzoW
xRcJdT8FLNfE8aSroVUUhSL1qbknja8wmGYsy9Es4NVUiUp1ovZJx1f+z29+582CiBMBvHoc+sPv
Ywtjh20A6Ue/sNM9o/Mju5vw6jo/s34rn5PKyBI6+L7IZCkqlWgeXToSW2haYLiXauYpjJF3pvON
+4teU/bpKTdPdwbcocPa4aN7kzO1OyrsN49ZmbI1VX/BX6RrPJqHfKT/1cRJwiVWU17mx19Cm1G6
qiT1yvsF2M1PRXhRftbSK69X5FxYNwReZbQvtkAR27ZM2iiY7ct8U7O1hxquxiei5tBfZpALnR7f
/uqqoPOlnDGSu7sRIp6qfM5oWvsOmrcU0wMWJcsKwfzbIV5kNuFh8n3dbumf0PoR3GWa4YsmEZX5
HM4q9JW/DWPPoXQrTrX4W6e8JKTsHO1BHPcfyABlghmmbtsVXgh6JqHDBiazgtTqLLe/f+o9vuep
k4fdyJeca/r2Hpesk6bMCRPh0HwFN4v5L8lWAW4el6ELshoTBcVNjsJ4CiIeME1q/fgjtC/QRePq
Va4kKmRcK64kyMRSieJo4e8XMkFrSzbMP1Z2mjJaIRr1MN5HRSYh/SdPD9HGlZutmCuvue/Q+xyP
jfUbQji+VmAjL0+WpkeMTK93kJ4Gbijg39aiuXQaRuXPr6TDdY8bC5tcC4SxqVBF8Rdr8umikwW6
z+5bVTo1CpTkyEYhbOpGriB9hm88DBZy9R4c9dq/8O2YvUgU6CogkAbHfti9a2QQKL2JCn8oVBTd
tfm8upMbIyL7W2MdwZRLN/wIXkGtDKwkyEFrISlBqy/MoXApQNuPQREaewg1ENtUGTIUG5ULx1bs
JgDw7bDGwM8Asr5NGSIv6L6pjXyPY41qF7jsALwma+dmykdIdLPC8ppRSXbP1Nc+xebRl8RydkFl
e9XyVSW+8I89oC4Hb2Ruaw/zGx/p3yBtfUzSN/9B6D3N50/ks2Ail+vFGgtFPtMODt5nzCAnLqam
R9/UktqQkRkZgzonBNRAUHuTNwCPEn6ItgycqMhpWzfzHtVvTTOxlFRgY/uEGNFLZdzReXseRCrC
g0FiV+WQ8+MVZZkqutM0aW4MjAnW/Hoy/iqe5TaJsqJG4QCDoZCvP1LMfmxs/Rl+0e8XcGLOqs6P
RCJIT0jwaYCxUSX6FqYxKy6bpYqpJd7aFwOE4Gbs/8V+wWHnldlxx0VcbMifH6Sjx5CH4HjGbDvd
J7yqP+bENke9MK0JZL2BmaLqJeFhbNZGwBNhhDc+aY9CTnLZG6FkSbP3KG91QvkxO/F6K+HHPlsJ
7I/AQKcryw1rLUzkTpIHj75nHzj/rLt7+6pJvNUDTV5pPg1IHIbYPJDDHGpToU55rGHMdeARDO5p
S7EFtYklCoiGJ3eK8cWD0gJeczQUtZxwwXjDDRPSkpIeaX3G0WP++nsm8vkZdPZ3LwB3A2cQqjHY
kkR9x4n3x+fysgWavbHwshM1NMRS9TD+/CG5BYsOlyZDLXNN46AMI7u9N4cG6LM3t50AScv2XMNI
ngZyZ0lxergJjdLfy4b0f7jM/vbfe7BavIWsVq9uxHqa32Hx9A7A1VgRWVpC3b86M1yJBsxkcon0
pPrAAeV1f72CkXQG0rNDffDiS74ovAPEQi9kVeySCwGBzuPAtqrfzw8TUfLPNZPQnymVbOZPDnU3
2o/qIbhVzgn8aQodYtyQxEcbVsIH8GhVujnM6ew5lHR6Mus+Jm7hRU2QGwLshw/Zifpnu02HJYtR
a9RHXB6VXB95reDAWAYcxEk3ciYpTITSwWBDRq03XJ2oBXFZ3wi5URVkX7l9NneqFGWTIT0QCjU/
x01uXtHhdN1ZQnN1RzXg7Z+8IVpCi66lmL8t09qoSIVK3bjWIfKopce7h98UPXTOlFPO6fzi7mpd
ReXKckU9Xqob8I0MCekxXhA1fuIlfQjRLEOMHlvA5bpeQaWsamwnt2JLdCgBwx47D5wAWV1tyO/F
E23BUUOV53H9ItknmdzzhzEwNQanME8rDbCeyb5V81uZ1Vgnev/xrf9Zbj57rgKojivdnWjbYIAI
G2ngmUtwolg1qowZMpOHcMnIt+BukzUzZXnN/WxczaPLuhUOkLfqdfOTRWsvRm8fxBvJq0hrmdFJ
pQEAeD0DDB7S2/YOHVMIVBT+lHJAIQLh7oZ0UiXq44IFOl1vrVK6AlG9zH8t2Qh59HJ3KtGpJ+yv
Zxfekht6NthZ0A01nu+i+I2u3mqZ4mHrz5hyKV/JqkWTSZDyXVF8kxAMSq9BYfDvk8VVjDg76EO4
iWYJKOMizg8K0O5g2/4pMiab1lZoooFrmwJ0nXCOjLSETzNe/82IM6n6Y7Wpl39c5nyHpxMG4p78
hsblHpKoTiP/10rLAZlk3F+sPeGBYliNUuJN4DHuKhOOpG7VGm276PcvyeXkCHtgqkKbHYVQ/wBo
sWzKp3YmqHGVlSFlJVs3R8EY64erqCQasZ5NfjOIpaQtzO4O3BsZjULdk8s5HSvHstKwEkfGtP7u
EtcSYFniCpjirgvU1pEa67GQFZcbmjyFiivTnOTCG/NqmsFXp2RBuheNYc9wVBiv0dNd2MXGgzh1
s3eDdTWVHhsLigfox2I+Yo4oKuyZJ+0NhcC45AEtC38JYrCDzH22AMZSeaOlHPL9/SdLqIdH2SFb
zNpKvR/m6+L/6YO2WNZhOeTMW8dCjcdQmfH94SEIrXJbXmSDgnZCYfDBV03bj2k2jez9bmFPwFli
pE1mTcf8WWXgvIAPpwfrCohp+eS6wlPc6LgUaLSO9LS5YgG1a9vGDdFQ5PjqiLT27auT+qxjU5Bj
RvSK6+e3+kwsvlWx8mK0XSQ3By9S3p+G2D502jPPY3CbsKwfx85MomGD07baH+bHX2uM6s1SltU9
/hf/5yKxVCFzvDy9F3/dOEARr0S63SvybtkYX6kShqftcNup3ERIpk1IwwOSn5yDjwYklvqkGNrG
uMwn+H4nMtk6+peltcDFYtrZ9ASD4qaRuxj8oyyJCThAYqExHYZAPNMInscYjm9+VeER0s2Zqi9V
b3lSUZ8dJRkxlESjuFwDrjDDfNlgeHoRzgOKTj0M4yJzQRHc5uYGv2ede/vOnAW1GXJA/4s+K/oN
DGxMq2g+xPmDrdxfX3k+iBAivrENlPtLtU6TJIn4iNgD+H2rbPSW0OR/YzRACrzXDKPjCnemZt5q
8kYEtoAHk/6EaalyWOQwQgjDORu9DWaoeJFnxgADziaraWTlXjXkQR5sJ1aaSf7dKvtI6TgY1F3i
s3d/1s+jO98tjPZPiHk+hwVkTgYfhgFYaEQ5fQYKcY6KeLcePMISGwSJawntReTIGulXfkWyys5V
mU+73eQ/NnwuO917nLQPylTmvvOZcKDSeMoEuxKdg1ecI6IBDoYZNE8ay8lI+D9HcUTvbJh3njtK
995tTg78Y0Sgzm2YU3Y4kRxBaZpxeFrp8euMcR9EpCsxzB7kX624AYCdE2+qn1BHN+CrPKT8LZ72
PCykWTQar0HHuNq37FQ9BdcHABsLaKQZmx2BvoP7BGyjAiD//7EafZO/wnrFkkPL87IQQoWzHu7Z
Ky9zkN/9Bb0yZN1vXpHG5ijDwDdawN+buebgYNNiamUqU+w9lW/kwkJYymYxBFAZNnaXKRTv8TkU
xgS5SWotdpK1G2+G0Lhe96LquyW4Xc4MevejhF4uhFkPb20m8uhAJv/KyDd9Q5Bhxl+MJgmf7N5V
E9d6bX6b+M/BSiFho5mJvDm+pPY67KJUEXlgd4yvimd9xbAzLf4IUFz78Z7A5okvNEjs4RdpSA6x
9kmGTxx2K1Y8R01qwsWA51V35Y+r+y2+zeHb/HczGullUD8yYZf2Mtf1svLdzGBNpVOy9TIZ/Ez6
HdycWMrlinfPHjA0OkYhQ6Yl8mC63wTiCu/tmyEWdL5pYI9Cd2r5DbAhcjS2K9n4KwlQfXnP2dJz
GxtBGGL4atDNdHI4jdxOxaag4+T0aPuEAKUiwq+XgX/s6/LpX6T9O//xBrr/avEfixKKGpQwjH7s
xLSdmkLNJJmubZ8ZyZHyj6EqRWUgAfUHFt5u70kobBr8FzNys4pyfZnxp6NhoidnPKzXYuXqyxJY
oePDl803cFy9WBgSL89rJNgj1EHQoD8XuNiIhqnsuvKhS3hkqbGrwppkR5+7mR1i8KO3jX8AMvYU
xOxr+0+/xCLzoMCUfiFFV73r9fu+FBWTP+futn9/wH7sG/nbB5AaTUTI9hC2zgc+4EC4OkFU9E4h
fhYREY0I5f8wXTj3EPcgnfThDxngNLCnTzDq8pCFC52ZVp97L5hyyGbOBIgDdwilXQ87U5yGFucP
+pBRJAESxZZsB7Nq2mQfdrqiu0iB+lNH5c/ShX+dz09530EG2VVic6dFwovMEjmvnGwvi7RuYMYo
CDkc9OcEKLN4Y9onTgMAOTNFDsYGZYOS07zijW+VS5tSuO27/NcAKx1vPryvrTM2kla9bS9HVMS3
FFaAB6MMZVJvJ6zxpIsDkb9ej5fPbXx53wNkvWZ0ob2RPfk6Wk9LXBg2ITrlkX4OiSn0XkWab1DR
MvGrQd6DyLCUKK+fqlYzYgLkaiDmQfYEnx3Rv90kbsIY4anMO10k9uapHtX0WhyrZJw//3iVvZb2
1QlqSSIExqHboHnDSbnISHCXIAuTwYsslTtwSJ3zU6LGuJSTG9gsg4itDaWWbIzqB7+vJBemAGHl
E0Q8R70EPRSd8op787ZsiV4leSdmeK9Y4KHm/Yjw+DcFFcRjVilykQ8DHESXKwPeHLdrfdEd6ObB
CXk2766KnYRrmhKGgjouq03YlzVrE4CD5ZNsYDy8dsNbs7xhEAIRauripYYm/55s2AxQnpRhaDrQ
RwdLNUF5fr5Czjqbr6glfAfMGdI98COqvzhxUBOS/CYAXl0x7qMssXrFdgTsKjySwss8+tEzfduX
FXTjeGyDqQ6SFiNdoHUe/QEbBUqstpYIV0sibLpJ0ZtyIHrs0GSlSU1hf2rxFlmQS85RnMa/z/Xa
cCDMGrH6W22x0J+2Ic8X3VlF3sk41KWnwxELrXUtDB/GaepBx2MjOAtsjnxXIsSIc+Tsuon/ylwQ
ye1h6ZKV9G9hAM6YHgNuo2E5Uqpb7kVfdG9q3aXgFnWlV6bFDHDgXOcL6KdJDwlJpNvqC73U8t1p
zBC1yTNQJlD88v5sPPAoUcWp3x7HZt7Bym2wTj0zeCO3pDGzx18GatiNyjZxJKlwZK+8Is0qB+2D
Ou74x2yqZl9xOCG7yZNuLJx0qlgpZuczaLRdRO9F+7BILF9cGfisPhpbNlrMeBZej7gXS4yFoEMn
Qia07EyTEspkQWl4NulLMTmsyX55peQmcZIGDi300QNCBWWJrU7/jaWrWCrtNeX8z7y9YH1W3ezr
EDhNfAcFJuFbSm/+fnrvIOO/dDmPMyp6FzS0Y20+VDZg4w+s9Q41+sb/yfMtecukeRAl9BBtRHPq
X2TG1QA4PPpHu6xAe3XiAtgmLkipJnuMDDM/Svx1utjKsWwbqsrxi3o8Rx1WNNBPwBNaVYUBfpXl
VqGUb881Cs3uShGthFYcrMT6ZH0ZYaFAAogiNx81UrHSfx/OJwOIcqk7P4JbxEDx3C+6QQ1mpDq9
fYcjKy3RQXUWXVyPVKd69uqsrX103UgU/vbha4TLvQSHIiDqOpnj+/VSAWRvA3ZFBFAVkDe+b6uw
rM6n5Pz/L6cHkgQomq4XlJHD8BdurLR6M0co4kE0FwUGogLwfJb0muf9olBq3pmp1DlW2rSKwWbA
5K+WMoC7HadNiibWzleRw1tqcN+EMfMZPdaorW6CNwUrEKIdMfzkkIcGxnNsxU0oVgXqfHbNNGaD
1ax/OUOyZoeD9RWmh6l9KG4+hQZ/wB2jvE9i3wZMKMiLOIgBsDxRey9JTbtjsSsqT45l/7DQVB0+
KSJXssXf02WGkbhIBwHIeJ0YT8AgLEwaU2/5udc9hVfPtkzgup4DKkuIaCgH69Rs8J3oJEeL7Bti
NDIehM5YiK2+KQXbxksxI/b0T8AGbXM9MPWYlW25448zCuHiB+siu8Fez0DAmkwNWvYbj8mKXsIZ
3VVNG7r+v6+Fw6I1qE2dgvwVpFh8cDiSRbFoH3K7VcTQLmA3k/a3w/39gfFyKs8YibAmqGbFAuFy
8t9kTbad3jucx5zFPIzfzMAQJVEQ1tScaVNrNB9z7yvnWl9Tcdho5WI1p9MpAceIXxf9CiUUFfCS
Khi7L9Cc4XNIU1OXvYBJSlKcV3pVEOTIPztoeVVv4Xal564PksaZrnajMNGCoo6WbJeJ33UaCXVM
4fxAL0XNTIutC0zws4vDXiyjH9/wUPpCouNmIm3P0fXKHGUwv+e8EKZ0cwg6YRlGKs9tizeg6jZ1
6kGTCnxOR3cnJiNHI8JkbVgmtG+Ra9xPXb8qysmXgqbCEcOOC+SwXWjgCGevyYhN3yTN1VIkZ2fg
p5kdTKXIQ1ffSX0MxPk2+oUrwswLKGlmutwIY2m6NloAvhwqj8NxHJpVQIB/IihquK+r3sWiNAaA
c77pIG6lSnwA9JeyjkqEPjN4n0as0Y1ECYJB9mUeHOQR7/dHUlrnbH92Q/7Ni12uivEKw0ynqlQw
+XUJl/sXkLwGkXiYQQA6DHqp47BQbsPmoPiiVhON2tDu+VSuh9pb/UNcMzdCWSck4N/qCBgKqSto
6flf4ZFYc18z75yz+psTZxblUWZ6WB9Cwu6gLudRGmZ9d3L+c8zTDsuJDf/YzaCygrrz4PdIuxtM
tCF0r9iisP3s4e2GAKv7P0RBIu+eNpezwW85O42HxFo3nbscOO9F6YSgQdr4lngIrzLs7+T5a+/J
6777XhYAXmnHPJA9fj1ntaN+JzsAwyTbKPkzshwu/XmOwidSzOMdSIGYPq6zi0wRHNHaUxw4Mlw2
dNr7VySTBHKFElj1AkvJO5G3QDxBd1A9Cz0+5czOwo4tf+x4MiiUx+PxOA0+FiSShAGy4xwT6ZlC
jBwClmunxD1Ca8lwi4/uabMEoaVM0GF+3UXAazlUX78PYjpuRbqSRFL67pINziKRXQtKAjTR4vJq
Py+pz4KtT0YPi0Cinh6VTIy+nERbPWzS0qhsuz3MHX5sep5A8d0iIXMTU17tsZaQdKTEOom2FErh
MlajP5yyOwGU6Fzb+iQa0p6o8VeTdIa7QMXC7pElOINY8Qxz0kdGOr/LInTRaED4JZ8O8Ojrj0V6
iBNA5kmZt2DmL2492ew7OmMvcOeEXXp94X9xpWzGjfTuAhPbJg7hcvA7ZZ3zngld5Ivwe4uhRO9w
Sg/FfyyYrn9iO0yiJB0CsgK0A4nH5GXne3hufI5PQS5dbmiwnpNkL/Wy+S7kdWIBpSfyOlYAwpIX
slrSNQIUnJP8t1ZdPo1qHc6zPc9XHDnfeWGBGBhF+HCxWAEWpsJ4MuWqupdIfDTXonn9YcoWBln8
PRBiKEdQEvcQq/KgayrfulKPn8gZu7kJM9OHKGUMB8sh48sUTlzxypn4BgN9LmPxoQKvz/qOLUX6
vZZdeD+za0fRGgbpras7TdoCEBfwghz4H59UbI5uXpobrnFs0l7qS1dG/cLwEtcA960RWjVDBcRF
WL+0j4HWOtYEFUDSICdgDQrXDss+f054DbPK5kj6TL7PF/uIrKu7IiiDt5eyHshUdzuXXZrHgvWQ
J6LWIEiUoCwXLh8LXg5i/M8mu/azp+W9VobWoNkt/WXjB7Y5Rw8e6HkWsmFk5DsXI3LKsTcj9jEJ
zU6VyTuiK59VIoygLONw3I4J/vJlpiu3UBdwzHHdZI/ZiIm9DeM3GeDP/bFaEG1TzFjAb0f5FO/9
wISsb545XdfE6Jb4bsx0MXhGFL038U5BOVy+n7cFp5TSWr0xneCLSH388aP8piPaC9AHdes3gick
ttGitUvQIxpvcQVH8QPPC+eM+hz4qfGECf14BS6ZeseTwULDEncgYLHoja7jGO1+KfzyrQJRn9UN
hA7E8EEpESlrbAgfLr7+zH6mlbztgo3VZoZF2WdTr2P6041+cAUP6ydGwqybDi2uwGxh+ygdWshh
R71H3NSEfaEdId2Isv211UFJ0jJuFHDmVYN86/yVPQEaUt6PP1Tvf4ydGRWZOpVQShLprxCwY4yO
opAlU3Gop40vqdr4SIfsjDC5MxTNTwhBof0oNJbTDd7UJTEXh17lNKd2uLb7Ff6cuiXQil8wu1wl
W33TUiJ9qyn2a9Ts6acDSdvBoOtS28zsMVgiO20g2lDWMJjSy5AdtZxOFoFh5+oHU6N/b24z7Lq5
S3DDirPIiSe6EOxBVKA/P+kbSug26OoCPjIsAhLHiTAGMERoKkYpOpnmcRF/pw0MSbHN3T8F+jV8
JafiCiThSaswds3m98opeXjGJyK1NjmRM9IvtfND7jvgh9O8gfR3Osxtt6EFCx5naRCqp6/mbGRc
H8Tl+HXDRc6v7pX/U7ybsxz83tArVVaIn1FhlwiX92GOFOWnpzcNiwXnDOLMluMBRZDGH0+wUuxX
0OknfvBR99aJsJ2s1uchmD6D54ytPRZRaVLEXs4qJBv3cxEyByAxeM2CvIWtQ7P3rXwuDQXUj6/I
9DtOtg63Di10yZUrZ/RjV/3n3S8NuYGerFwM1dE71Q4VNsjMU8gcpoRn/zDe8QZpCtK5tWF1IXoo
3026xso+9nnXYHcuC27xg97S+2hV1eReuFVx/Fvw0Ag9WXU+5AXKzK5U3RyD7ERfrcHks9K3Jsc2
9NCTZaWwlybAhvzUjpF1aa9Cu0a9UIFWsBrqkRripDXLe+sqfz7V2nm7jFhwlLPdR/Xt9hHhT0qr
LPhCDao/HbISz4QiP+xmxr/RJJpohV5MTmiW+XRFYDvJnZoxfTpHDEAgId214IDsI1nClfbshPev
Snx/sv9qbl1/cZpRF5yf/JGZISS0idQMcqcZuUuTOzWX6KYOP55DW3Jz/pzX4VE7mkrFQh35Ol/1
jQwI6K4fRwkmcl3vkDZZ/mzRUK6fZnw4eLhzHXDcPCedtXyOvErCvGrj7d+K2tOf+80fP3P3yWZ7
j5PXZCmqCwj20yJbWXQdliPgXQGUAnNAWl6x2OiFLtjeNpsT7dI7bouC5ZMnGjJBy+r13RTC5Y6o
XAM3GxumGuE59hr7fZJy1Rlp5+5BQgn0xdtBXMUWj05BKkQfwXuav7UqPEpoyLGr7pzGeVWk2ywG
K2qZJa1Pi8lFDmFD0y5ueSf77q0rJgJwpEVivqhZXVIFTt0ike7Ov7ZTTPJth4DMtHr6IdkP5hv/
8x/83cNrT4nKZjSSx5/M22/ILARUfuqZruMuSHuO21gGXut8QhTx/kkQmOxUVv+jaV0k9qL+gCaL
AjR8EF29EigV7CR0vEzENstZjI+5kv+pSMbzZiDRe3XKnJSq6JGtV3BUTHCXV/dG5vr1mOqLHVPc
UiKFFGu4Ii7yEm+mxjazV9PTfgxXkHJW+TPZS56TT0ydfvZKPdy6XfVS4eDK/3hgk7yBB//CP+5y
WPY4XE/mEYBOkWc8vP5PnMPTN2pzfovrYmpZAqWD0CzdQuQ/mJWJaxJkHt161TK1L8pkgOCi6MwH
qV11VEnk9AhNy7ROkiv+E8pIAriRhMJQBouT39WUVGBo9lHIRaBiBttUhfAiA8ICTU2ls+eaZOKC
jqqy4NeW2jYZVgGwpD3VSsk87ycDNHo4+q2/XfNFJU86NWh6XvS0SssczCBDyLsw2EpcX0ogBB2V
TbucfX+FTUI895GBRG9q5w3b6PLrf6kE3XPoujIL9OOmKOkCsaq1zrNs0KxujrhOMCKHxmHYCc06
/XPZynGiGwCKcwXnENhLJx8x7vgwDLJOKHuZieCssps8ZWjCJHhcEdQkAXXx57TN2tx/9NeoHTqW
YUHju6zFYhXI3LC0JGYFYAdUQNwAzpQXfH0EUuIk9e1Pw5T9PH6N5WhBeEnvxzthh7K5lju16YDb
B16jAJIzqPOaqbuWCeeMPFzjJaAkJiO1haEbH1jXlTQLgHGS2TlaTbTpxNap6WEQBK6gL4BZd754
fDIvUl9uYtWlZIj7CxWeYG27yvG8ikOB+HJklKIFnwqJmF21bAoN0jTFdTAEJs8yVKiXvSkZSVEe
/9MIm6kZIFlRQhHbE/NYkgpJsDcGTYHq9XACPt6QQbdmgsPzZFAshCnzanjrT5nAjFHsjTwxRh8O
8WbZkw27sMQV7UBeG4TOta4z+uXabrFT8iXuiOXni0Lao9WWvjUVn6r8HapGHChGHFB9LfHZeHFy
HaYa2c3TCy7gryEQXcn9Z2MDgFuliOzaqnGXSOFfH+fGTKnPPfkvYsn2UN7H0COpqyEpohFDhyE0
kYADNnwmJvJ1Q9g8ve11vh++sk56A06R3DvHrPyixX4WzcUh32E0nMKQNN1DsWyborQadGxJniNq
r890Nnqs90ReHvrHR9N9o/PAyXkv+lqvi9aK99XkNg/335GP8qRiT9+l1D+CKtFJyojMPtbI0PKu
vBgv7J7PaSc9Kgzd5SJNMraBTdTOyYxrTL8qLQH8QnGz5a607JmA826q45h1Lm5vSZDLRc8yzwfZ
xpMh7rLalOnGv5w+fs1OvGDrPj39p7WK9zKMTMBqf1w1WG9qngc6r5l41K+ABJeuVE3KozmOFtCQ
7NnUsjVhJOzRUbI8NPG8KZ/B9iaYSYLGiZ3Je3c87ukdkBLgUy+fLOu411jXAl43WnM76FxjvoHQ
EBmvK5BPIhRaIS/BjiHnfalwFurBw+GXfT2kTsTHP52gEPD8xFjNymYCVqiJBsKCjczyLG0/kdO6
TCj2dKRVZMwkTYwvHfCOUxJwfgeUuD9MoPfl9JCFvCglaH/L541HqgjLMhoS1WL/E2wG+dS4wMU0
AupVYuPVwXfM+Af2rQA9nXBH4nJa+LgWIw5Bh3P1ZOmCNwM/PO9iCtIc3DsxQNWbtVjod+pkfpxX
MHiC7jUpe4+gAhAGckarXFAfQF5gXRGyl8XQToOx/0iOA2uL7YGUE/O1Q+xkYnd86oOpEBPymT0l
C5lJz21g8zjKiiojkHboCywge2QMtHdFRgJbSKnQoPzDEzimi47oqBs5mnyWD2usbCtCQmdXmLcw
ZyUz1m37rWWuaEQTjWm0eKb7nFPPYkiRY2rXokhxQpwZaPnkgR4uujExKtjWQAQcNY1B1rd/Awdm
Ie1waQCKEc3pGcchFR2bq+SKenH1gO8lCSvLU1svXg9y2PDb2Zz+NmBzUw8Hc5XD/O5QDlAafOhz
oo+aAqvvKi1oRmQdgaFUqlS7KPmLSuoow5ScZmXu+avuSIFqoQ7bBFdiou3ewMeIymVuRL5NZMWH
jetKLy0Alkm8O8OKv3E7HqbF+E0OnAHuLsr6y6vx7N9NXUZAYEBNm2eUpBBOU6qxNiN2SQ+dOUdS
bRnenMRJ4nflsbm/RZsQLoJU97HDyKduWeqZNDAurLfaG+bsGPv9Mj7EpLBvCwTSfCPN3RBAxfr1
IjxUFKZ7Chfp0W1n7H+JZF7zQsBaMLPSjPfVncxW/CEQBykgth1Dw67ANjveWgkVgb4b7b2Rzncv
IJ7zSnA5RnsBOsvOVuuuzedVOBwZPGYi5v+pwOATjzgowNHmM9OqtPlcUm5MuU4npytk/HqwAHxW
+bacKma3L/BH8UyIzxeMt1ks7FaxpgPAOJfGa+vMeRVN62nYQOV8GfraNwd6OfGF/LWwcyTMaynw
PitaZSf5ZgtX9okhL+86GuihBQwsxPPkGOM8JD7EWolK5pCFa2W2jG5LOxJo7TFazWjU5q79vG0C
eye2Y9HnKrddAThOYyUJ8GIoCOICROwME6dwJtY7pR1D8WrtrPBVXyiK6/H+xE7ceNWzwyF+87QA
eJf7gF8IVbm5KM++w+tWozDlCiKSSBm5rYpIJhCk9XasogvhmcP9kvNaOU0nPM2ZwASp57ZgdDJI
4WwVnHHdmNiAe/nmly/YTWjqjjuGp9KYnP+wAuN9mCga2OIJnRn5BiCFlSRyhDbDGdCUlGdUFZL4
zetzShfEW+sFGoBYkLbVU0vOnfcYPh3BhEfvPGGnd71EqYe3OWvdlOPA+OWy1TDdrZ0oeH57F3BK
Gva/QV0RVdzBDbATPS0BahqVhTUfb2FbEPCZTdWO6mK39VX32eXnb2qs8z6B9wYHpEsPh76LsYP0
asQk/Xtge4NPpudbsvKvq7bvSIIe2Rqb/TZvBobI7mk8I64x2VladY1j1gtgobXrusvn/Nn1dvei
9590EI7IQMKEjaXha8m5iMQ6qUCvZuwFbBVEhLDfbdlyzlbNwdnGGSTkvjaUPT6jBVn0tc3Rro7q
3tlC7anpB2ARt6hgjgz8Ta5bPqdS9R1UOb4psS8LXe++bZykCgw1SqgKR363flI58WteRGY83xk9
dnOhr915WiC51Ch5qvH9nNevSSyiagu4QclPMo3hbMcepKVs1jG8gT4aJg660WvU9uHQFQHYn6p2
OQ3ye/Sc2u95jTjRtG3QKY6P8ZX8FUG0afO7sqVFyKC0PzKXk8AnIV/yOlbbIzFcgWCPSwUv/LXd
bNmnhroxgER0CMO9vyvDVoyQ0aCBtKK4NTKF4UBm7vA8W229BBsD4HM91zKPueFEKLUz3uIEiTBf
Xvkj2//+AKM9wUV3ltKtG/clGINL1627l1gTNjOpqg6MtremVoSU83dx94oRJXOkfX+JtSEIj6XJ
w7MYRTjFTekiRFNy0szD5lmKn5xTBMtkJwbD7E0virsb14Xqhwt/j22RszHjzT6V11p+MZqp5IuF
ZP9ooUVtmlho+MMetvMQwJlbouDJRNlVeuyZX5gL4thPz/VR9SamSBI0ohKoBcK+V8AAvgX3qMMe
xRA9K7T/YgVDrLBjtEIK7trPzIpr+0qrkxDeHbI9J0H5XAgjPgMbCQM+TfnFT70UeUVaKfupnjep
hI9Kwjkpklu/Pd2Q5PLwXbjilhsQBiOsvbyjfEGVZuP7cj3/vddcrAdsXr9bRzhm2Fs+xp9/akIu
xxPCsliZWDkDhcOvLgcY5FNfZjT7+bL9UggJzRZ92jrOg+40n+/Pcv3FVNWVkBOEDoZJ579wwbCM
QS0suRIHPNUQBxeNco7LYALPfLUG4y710Vg23/wq/DxkEXQjXQl9FkSVmHNrJzEEbsdWC9DhIxh/
Crp3zaC9sq8bor0+ziCXMA/BNi28GsRZ1e9SMTm7MqJSW56UINeb3Ul9oC8Zvd8VjVs/uSoPJJSo
wde2MdyY+8zMx0rg7sM+cjrvi4jiEpMRvNdz4yyS/tpmK6F9p1D8dl2eRybda1EUIB7cOnP3W5/o
fGgggXuIGX9yXGvd/1lvp9qS7oiYA2aSa9NJ4OQObiWxdOZ0ciXDpWOKSlynMq/A/j0RTCl9fCMV
QGqA5Gcs2MyIswtPDCk3vGOmC0xpm+IMRvWXXP4Z15eqSt0+FBvahm7HFfRzbN8GV+hpQnnHxhnb
vEUzZLyFawWrMz8AF0onpBt1AAugRYwDyh92l9BOFnqqLyRCsA3hE3ZkovZUwAyRRpQbXJunvb3k
6r5JgBkU3LX+dkAWKrdWfjYrPvgf3wxKjHFn9wTFjgoIlQg12Ar0mal2E5az2lGX/knBrQpEmKxw
Xo23bZm49dU48QarMr9ExHFb5mKdAv9chxYyo0/wowIUmUmcvgSMKWYIeGCFVVxiKuYIhsK3gMCQ
5HmCtMP+XhWyIm3wK3jbqDBJbeon+YwozzUTSbKjAh6iSKxFwOjMCNa25IW76HLV0An9EqF7JY9K
uihb3gsRPuN4CmsdsJ4thrlXsm+MyDMqJ8pUm7kv/B2A9sANALCUm7EdVph5ZKgE9bssUm1I6sj7
0aAq4ztWAKN5/a4YG3yPA43MqlzDPANtH4LNUy3piiShldqsV8ycKD+LTpE/nrRYsZHO8WH6MmiL
hQEXMHaQxlSuZtRqX+9aplXC85xilq0sxImwBpa2l3cKCeIbexTsY1pMu8JwctM3pgMKCVQnk9Fo
yqKbOh1yYC8kVpiBp2mz2WHoRQB3hsyEE2jzixG6tSKREqgv1BGN45srUtAYnGz0SKZla10sN22M
Ulr2ixFwirpATktczhoQOqh3jXjloLIv4ina0Yx8rCI/qe6jssmwi0EPXrICmSWmnWwtPAkJG98V
pSfnz3jrFUJAKU/VTtDPUCICZrY+0/VeW056dLo/kGZydovqofF+/GL5asV2C7ieY83pozbkKF1T
vrdU6HYXijCfqoyHiv7ZeVJ5YRySYJAe4Dcq10aKoCKUqWKiTBIL5R1dZThVJSKk6dHg6gtPhtyT
ohYd71Xk2jOx1MfdQUXOJgsFmyhUMPUihkvNmI4DaE7cWbP98i/vV4czuxi5qNq0Cv6Kbsk/Cv6n
4VsnZtgkwRfUjtFg4hTQeJtJSlCtIoJXCEyoqY7micOT/vwisEO9tgbdTi0xdqgkJ1OKeZnB14b5
nOwdmfNrwJf+IlAGfrCuQqubLEOljbGe+ebRaesWjs7KGE9vqsPRFnI1mrVLERJiugXrMa0XU8Jl
T1bW629nPjbku/d9R3ncXJ9fw+uCetBfFCsZ057ygxn3fSprz5JL4AOUWtfkXXNyhpxHYmMU4WYN
bWdHwyFHYanZx6vXXYrNUaXSoPx4N66zSuJzodt7qVkUvRdFhrhELB4BQGWiU5JPg0JvjqMUYEds
bF14E2/ZTBiE7/kss1PzHjWGJ3OnfPVJOunbiu9Y8khIQSNP2R/c3AwHZNYQIyDEoKcQ1Ikgo2Fp
WUPztVKnQFXAC5pb0iq/6HgSif7vSJnQ9lvSasXLO/nuPW2wB8M0teOFvQzv0s6I40OgSkjWpDm1
shz0a+eZEDD4r2k8rt8weCllnxtVvOyIyYt668aKlk6DeSjBcdDFuQ1TGAdmhm010PrGx559s0Cy
2EevFA2co5SbUUSiQn0qUK+Wx+JHxAjlxDo1qt2DcL3GDbK69Rdj05GivJ8z6T9ecKTmT7lcAEA4
9nA03sBjVfGHHMpFav9UgSgpf9v36SC6AnmZ64qGDzN3Ryjic1bqmXJtn8Zcgz6fk9Izme0rRwGx
4qnvvIt+O1YrO24nIYNE9zgsICGcMOdNro11KbLpJpNQNcyqk8Nc2l66FmXOUR6SrN4ULOFcrhE3
k1Dr+GkxU6hRxgMSovRqdTBNFcmyGkJPkge1ZOhh3JHwi5izQAT6uetyPJpcsOsTlo4TSUHJugn4
JmvIrgUFL+jOGYu8Q/9FYOg3NmYnvWgjbvPKa/Fb+ePjdixGGyJ/moQ9/lop5Nw0Zt+sfkMtHvBa
PRtRvMLBFUz39zoGEnDo1fM+0tzHq6jSFYF4pf5p19woLhd9pJweJ4LKXG2f1XGAAvAOqc00NP2L
KC8i4yKoowKBNwgnvs/I7sUw5F1TJW6MgaAdKpBOYQH6AM1e3xYZHs2kaNH2E9XgE5+tGpGgSApA
H9jmfUxe1bSkshd4GvOsd7+IA+OK5/sitW9/9vyzm7YmcmETNilNDwU29J4zexzyiUyXt2kjfwFV
BFRcWbaO5VrqFNdKEj95RFLRJem2acyNGDfiJ+crpvHB9cT24kTzkzK+t3MgllQ5Fb1+scL4VwDO
BrtIKOt86tjc7heP/rqmvghIJGg9IBKMwQNkNrmQa4dVorqkQplR+IASAIuOmMJ2AaHrsUV3iwLY
budTo2UxyjSftByteyajvyiDbWH1yDPRzrLHEIHkZfKB8ja1TW8hyu7snlkl+NUBhc00TxlKT1O5
pTBmBizlEyhtNekNu0sQERWKGEROzlS789N89pCOjsiU4gF55OQj/bZ1LKp6T7zMJ6jxFBZDnOT3
saBFkQBU+qukw85+nzoXj6188NKJAbQYJQXs5DoeRdpfNb3hhUjiOtGMnVHkYCvNYj3c/hcg+3AW
KJqr2CVVVYOPNZz4CbYVnS8M11VijNVLzxgZfqUrzKV8pqg49PSbsyab4XYHrH4n3Ciibryagcyj
e/fyVhINlSd4lT15+I1K0Xej7l2U38QAnj2heXfv/upI3KYNWLaLBT2rquTcGeTe0IxZbG88hhvU
wgZhTi+L7CmrBV99U2sEZavX6d8xo5DCf4+9aeTbtI8s31Wy3iJe0EuUTuyLFMzFvex4jbKVErza
t4j0/mCjAwrztl6Bdmm0LxGWv4s/smI0LsXpHdGPU9oqRsnOyFa6aqG6e1ohG6ujpsLc3okgTgjf
g6Ec7JXT4fXSFdz2ELOnCbYt0Q2hM+41dnJ+cPCBclFZxRjTEaV7WqUbcKTW9/zg3zmgYIHcXqlR
zEgI/vvZF1HxbhPe1oegO/gWEbBIuP7rt7Am5H6XGPCyy7GQ/VSsUoBe4aaraD/57ed5bXQmKqqE
SCWXcdQKOzjVZJLpdtsRxal27QoxTSP4BhO+MsNu35d2P9nK5xfmraKntHlBQd5t4DytbVMePIaG
8JKEmTSxMMMC3IWz/TBEdvre3FumgAHyMHdL0dwkRnOWoDRhTF4MoeRrX3FUEK/8ZZz1KcjhVPgY
0Aev7GmwS3/kS7pHUfPPaM2JushU2K51Cb5wduDDuIcws3MCnGz3lztPtoGyqIOcFBPlwMsKyqQ5
EhT0XWYyLj7k2a4cbMzBUKr9/GjIbpRXJTaAuRT30YMI8/vHcRfWywRgq6Sa8Y+kwB93t2YKN7E7
P1uQ9pets+6n/6yK8y+wdN4Ts2moy6AANJoZxKZrI8A5xF0dtC+T57E3rng9zyR2YMa4huu3bi9q
Y17pzN2HVUzyzxMzjOBeYQMKTr5oCJkEYYNkxq8SIk8mmGXQ+5eR1a93yQv+6qBeHoPIcYO7++cQ
2yGCynd/+DNC9mIzcubAHZyKu7uV3VkpnFcyDA6Bgh1IXxzbvLiNO9e26WXBvB4J3D2yTyuoGvlq
c2hTyTeNwBUJvIC/qlDH9XeL9VKUTyFiOBwgTOzjUS8G0nGAQe59hQxT6B+ZoRABPdv39DQZFUI8
GhAFfltuEQygYwGVBzQk0A+lLhI29Jk88HfQUHKxPv7cdf20ejpml/SpYi7qd52drtEu1i5DXyGP
9UdgXmer0XZ5sAHtNp9hrepsH+UWdCGt5Jg8ZKTSNqhvg4smlsYJVNfAoFXRYPjmcNCUPT7+cAzX
AyANd4/qmG6H3syJ6FJ76ZTsjqzWFRZEPL3ZpbAI1CATNApldnelWgU1AoC8XS6FIiS+9dkesvkH
tnmvKXMusa8TvrV80WBYndxm/wF9oHmoobiBRKQjN45Sg6TQcwDk1b8beYlXtNUFj19vD3YeVWxl
/kbhlMp4YvPFiVc2LI5ozElMOI4RZlq+ktNemIY8wwFMHvsLejU2fkbFA7Zjk7veN6gIx9ILUJY1
KRTH7EH0bJ8QFeG7ebuObpjn01nylTZWNlcm9nDn4okkJja6OGihjSlNQ0GIbo6xk3gK1XtWmiUD
0w4m3xkJzVTrgQlHNNzd9n/hdqXDzr8/flBfRkbWJo9yzob7+36mnciom9xyVSeFNkoT94fj9Je8
ZGItviu+2fF3xH/47r4S3u3K0NP8I/+LOPFxI53LlG4pajcc0KwWvkq39varHv/Kxfp66Xpi7Q9+
AiB7QZNpDCb0cmbc1EwfjDQ5NWdhHvIypIwxtLLOvpdw9qM2ChyT9EaV+bUIKGFdUeUFY3CCPvYc
Nh9+m5Qj3rMc9OQY2uU9GjyuWUKjGsUQ/IYloyLaxFPKUijv7+Kb3rQwm/xC5iXVZDExOHa17Jbx
gZNgCD8P3HEuTE3ZSusCG1H88BesstSIm9MvXUX6CpwEVry5PoEgIDmU7MVHRRMX+oX8gdeWI/4I
rE3ErBtao0W3FgeGUDLF6UxAmYMVD4WR+CaWpEWsGbeEWrNpguD9lVE6JlV2TtxyzAcNMDbutSbl
hQcCGltFgnjRCGYV00rp/dbeTLENBuF+Tmrl6d7g89GMkrySuwhNVn1NKniVvJ2LCHenM6qe3XB4
5b00ANNFEP7tCX9TmRUjEY+heSsA0rez2mcqVqLCpxECH+F7G8ka0mqPEhkwqM5Lo4o2C/S+xq9X
XtoWpPE65vU8VjByU8x+Xx2IO6dlW1CfEwdA0YLHdhv5AMR/uchfI+RaJPcGMXY/xcIQ18Y9Z1to
SDqajxu3RtJpT5SLLekNaBzWNnRl+/4v0RNIk0c9h3l1d59ZeRPZINaK6Nw9tks40iS3av+hY7K+
vErjXZUKdD+8IHvVoyhy9Np79PD5RjP6TGK+6MYmuWTdcKo1cczX5mepdLjCvneq4ExO5RJMKY99
uL6qbdSC6r3qV9mRHMK0KDUEbAESWwTXtsDJ6xsUGKtDJggiDEr+NZwpOitTGp77LxwoUfcqGwtx
WVyff/HSyGC2BxCrU59Gr6OGUlmfmQnLL2Bt9eRIv/yUrPhi101t3waEUOVwb+gPbwfN7ZY9iNHZ
AVHFHtVGetYb9B+GpZbgJ3usgaexATgNMsgSu1hp7CT3Rl6R3EeuLnK+M0oJbm8CyTKvaXgu0mZw
FWI+l/tMOQEgx57I7C08cEMKIk13ELeNY+sDeU8v9lQqn4qPhy3W1i65gu+UYBnKwVszMmHnU9gD
ZVRe83lQaJJtcUcD78uIza0E/RO2NlYUoAfwc7ZFFMuQPplMiOsiQofq54Gwtj+IDUF3fcA/kd7h
tK80kqDhOIpUJ5qg1zwYfSItzYBE61A/H/ND7qvlXYR3yslpgpAkL/IW1tTnAv6rhVs44sv3Qv67
k8uSQU4y+dbP7dtBiGx0bxKiMW/Cj4D4eH9xyrT4diE8Lh99dc7JEO7BJZN4KfnTPrEp2NrYTKRa
EAO24JHI4PyQ4KZg01M21/CvGJQU1HIjTBiJ4rLlbOZcOpSSjWIk+Fj+IulskAS130pZbvLr1ASu
kDIwK983bYfa1/faYEAI5YmYfZ7rpScb4lrmhH7Nxvr4aFO/YKRtxmIyGmV05HPKmo8S2NDHwMwq
YS3LT/eGFpVyxqR+d5PHygl/kZvS6JntIpADkq2NZbslLjfiLO6H0mehacsqDCa6+nRVUKYbSE9e
1CAd112KD2dQ8zvmU8FEUuoMuJs8Pe1A+Tu87NljFJpuK22i2DQAlD5am2VwQ0VKV7+NeygBNv9u
r8qd9qQ6hDJ32Wo6SWCByNX6HkxkyWnAiZrtYjPufjS/cKgMprY/7mBklTyzZJs9iCaZJc+MnjiH
juNE7hM9ffOGnJ0EWX32V8zjljH+Il/h6NS7PnRssUyXaLwsLozShV+WJcI0VKvxafOBKj+F1XhT
LJcnvJcU/vGHoD8h2BAvnNKa5+/m2oRo41Wgs3MM6xOj0UA+7X5RgB4YBmaZYxNYxgACxIr/FPM6
YsPCLG2aJoM2Dz0yz/UaraWLEKS7KaOIFYTiviv8yKE+keO59EKHyjUkNODEpAC4qZK6iDYo+qLr
ZTh412Qght7a6HqMC3qo8Pt3TUhr0EC0SKKCLe0eLRHS2p3OoqDzEgPQQJJ409qZSSvz9eGslN8T
9XklhWs2Yonexb7iv7Mr1KQAHl1BMJxuSlrtLvlmNKdD3lYdkStDj+/e9ltgmFCJIEck4zL649SB
zqdBy9Y+p0MOAObPPCGBrjX/FBa3BIjJHWlZXJH5e9K6HDB65354uXKtBUy2bXvKgpeMN9smg0xb
2CBqVVHmcHANBLuuWmrFNof2mp5S2gGkCRotvIMGs9jdaW+0leRAzTUtq61xvPKwwkoO5hqL33Kl
u6mMSevXABRZ4hKlJRX97s5tereTe6TtPpHPNDA8CgGEee/EUp0C4gxj1NlVCdL3jByn5TFxg0Qs
uwJ3RjYgo2IFnYWlp93F6xxOCO5hqeKvYvDE3Mw2ZdF5JmsRZ763whvR3Fj+VAGp4Sm4TFKpP4K+
2ueOl4ppokxVh5LEBg8CIIj/5Fs6fidQoETvh52NWRT/Ji9YqLHgursnyNN2sqp3rHK8iAn4gLGX
Typp7qVCIB5muojkGxQXhwkAdcBEnt2CXemzw7rLaEMV7haOEiyaa5U2eyQGr3GmzEWqHhkSpLeB
UYWJWfq0LarpJF9ua27jijtD8AwHTi6B2Pio+cKuA25zm7NjQqHAwafvv38HieO2BSFE9wWf4ELv
MO3WcLQi29eeRZY031AcqzxP2Zmsda65t777htbwVumIQ7lIDs30YsPXVjbBYA/SLTDsJbLgHJPg
IliG1p4zUF8crB6ONeaOYKbPhs3BohRdNzZZo+oqUj7McPn7XgjiYAL3lMwzVZKo6Rhsp//DYQxX
71kZA9PSlSpqOUJqQGTLDl5F9okt8OU1Ynwc/0LPYux+UHEPrjp8/EvZGja2qdP69rRw7/RUoTeW
wSPFKTNZ8ri9zMDQf+cq1B4LvY/4lkxYAnUKInG9HkLsdnD1x59R5p6AyKeKrr4s8E6vUGM65WPO
YFtbGnilvtIp2fD3M3HKy35Va1zkVJInHonoKcfeVe8IyLl/R8W1Sro6M0/K7qICaWP/iPQUzTzO
9wFjPhULITuynzWdts/i2ip6GLXy+1BFZAmnH8p9oO4iJrEbgZIHfw582jBTeUnsf2r00WKoYQ3t
E9A1Rt5Nq6xcRnN6HS9S6WRToAQ2r/YZV8NRbincxBgc5WI76TejFp8CWQ8aMHTGieImpI8y5AAF
JJCKVOeOBCSrS8FrL5YgHObMvG4D1h0222t4v/4FGMqMuMWXbNpLodRR71NjWOxhE7QYdPIXRaPf
B3SQvpjVLBGk1jP41yT9KjnVNdoI/b+GtRooaHAfF37kyfvql3j1xM+vZSsUA8lLE52qVy1jhhPu
0KczAZa4Tke4QfmRiJV5tGNq84mBrZbGiHT4IXhlb0Qs+iyj9xEbx6La220S6puXek0Ob/Bskm37
pBZyW0hBBAsQ6QoXPe2SXaMyY1AMcmbMmPD0ENEiYFQr7Bo+pZBFWp+++3I+0nUbyDmGrZDd1+1Y
XfCUBD65/CSoYG2StD2WikTipABpM60Y8bf//IxUrYxaTPIuzPTaoo4Oq7xF0cZx9vLTosYjdYp0
MiuFHfc3NupY/lLQBZ8w3SmIwGtGFDDIv/uIWSc1F/9yiBRJbF+64hDEdsJSHNYSgyIKwkG1EoQU
C3KJwvhc+XvVreuBSfDSPuMb+ebYGlpZjXwvS2zPqSwdS0AJQ4cCBjdfSjMCc/D+qqaQlBkJ7GXJ
h4L0czJLw3jPiKWytXsQw6pfwB3bOqUDjsH7mUkrfYgPGV4JVb/gC6UAKdSS7XdAMPr/hiYagmyN
3GGvzvvTAsHpuI5OOHwYDQocxLacLK5iMUuSwQbYxK5y9Icyd1l0n/CI6UuxVd5Buj8gAAdZJ0gs
vsdk+VHjVupuGRJdNd0xPW2u/HT6cIKyGzu86BxsXUxF+iO9euLcP3YHYW6+FgNTcUiuhsRInMGt
GFgXfBuayWmB2uxfZur9LZ14H1U3LALe2B6JVgV5v1a524mI7UssLALMfa4iPk4Xe2Gzw6Cbd8/R
d7dDBROEJCXSMzSrOVts18XzZGNuQnvwa/mWRWyUZ6dLBA7A+qbSIoErSZblH7euy6YJ1Tvw5gIi
fXTSzQfAN73PGz9k7sxmxV8BHdd3ythFHdt0JElQ+AVw1H1kwbjPi31VyWy3VG7SIVyhqzLQPElq
C7CxFnyuvfMWtL43m0S98rUIYNWiV0jq2WkRb9NsPW0o9u5s7at871YWVUjAdX5mxiblQpsen5i7
KNJmu2hKBw40n8wjTwCVamhDyF3TGcYtwP5AuskQ+LO6UgGMNlGarO6PsblexAPn7rB1kaCizl3I
tWNai8S/QuS7TSmBpaMT3AfWJMcrqYFIt+TrY/3rmXBwSLbVMGp7q7rMGCyRu5JQtbaotc9SFb9Y
eP3Lk5oa2OKUuuN9reUkEWkzq+g9BrLcTagmF6MyjqoaV6KF45LPuq9C60HXZN7eu5kGxLFY4iFD
Sfa8pNOP220ho/7D99BGkIdY1thD57DJeKXBupK3ps8qwFEK6MGpO/CptrWwnDOAxZi/W97AA8B2
K+la8aEaWmvCdrEIm2cJ0JF2J5kUf3h7zzU09sUhzbXcQP2tHYmcSRagvgZCMbFX8IQHR0F7wdpi
xrAuLNncD5ipB6KMhXJd3szSHw5kDEf7LUGqNcqthgxfYv0avyP/DiqSHIycgl6xwvuzjOGRdX4R
YRKtnaC2uL/2Uh5hKuN4d4thLJ02naysy5tWaSU95qfBP2lm8Whs1JR+uvOOAcTQOI1gxnDN6fnX
pCchE2bWxeuj4d640Nzr7urA5rkeg41Algw2OcLo7HlUMmlc/E96QnEvaXjCnx4Bq6PwVmxS9XGV
yORV2AbI0pUhAEsFMOiiekCSlLWQ3rIBXxxdVdVUktPwYjeXJUphROrBb+5HFo7fYDQFNwealAAb
UwJUetVhUKrRem+DcDtioFlbt2JZHDL0c7dPAfZhXSnebMGL7IGC+kQwJbMlznsbdIvnSPnK774S
kPBBF8iMyTYfkJYQ1/CouLenv1j0EbFYy+CEW9Wnx7kh2vbqkWKtuVZpbCi20oR1ekQrk0081466
018+cYjzSO/lK0Nn8BbLZ4DK66NL8hrY1/7WU0hjyVVfesM6udRYoUqVLw8Ss+gzjdCSJETaY/Sp
yzeg97sTA9gA+gVYnDS6/OT/LxNHom6TybY3X7PWCnxrQEhu8BhI22vSGX+ZCoTiaX6nIgcHi2wA
FZsfPEdbVf4cfLHfyLAOszhiTxLYFubvSo0n0CN4TSuu3B6IscLLB+bj0/coNLeAabhH//5y4Prl
gEe8FfFm//vtPNkx6hegAxECp7rDpdy8ONeTEw7ObHN5TBFOTEF3lcWNydu6kFnUMts3VXxcMKza
gee1aYHPst6vGp4+VcRIOtdaT67QjTlI3ZBEkJsoeUOqLnBGlSeUQCucXlf4Y+0nOpconR9MrGma
sAztKK7xlvMLFYSAWlhegfblOyoz2T2dk/K6lJ7/YrBmV99YZdt68dNpilzAud1ENEJP1aX8Gvlb
IQ2GCiBQekBAif4JpnNH8ccSbrHdHjvdOR+inJGgi9rETw1QlzdOH8O4+feQEksRNpqfMkWYC7mR
gy2zmr34hoSMYmHpugSYYpahZklHcXyvOzBlRf5xkoHhXGayGLYkkB/a1F+IK3g0tUYDv9h/sDMU
CLN5/7MUmS+ttGE6ndH0wFNPcoN5aM/qaCwsIOwX1NMx671NRY2LRnbqjZWenZVDSF5lO/OZWMuP
i/8uqKD5r0mEhwWhF2IWD/uEITMIKqSVaH5NxxqVzf19aOzogyI0raFjeHLqBvaZ21T+LODMZkri
VgztX9XK7sETGUFFsf9HHP+Wtx3ZwoaBtlEHCro7Xmj28O4Kezq3UsfzQIOGcjNFxaOpm7s4llPU
DJce88sr83VIBILgw2EgjEMRI/C1OQqH92FFiutcRh7qOQmqmiPkQ6/cVUMl02CYtJhe2i3hfp+v
HcV9l7miKvXtyrmWIwZIG8NRTbE8CXanzArX+utP894oTctGaP0nZPawVha7ahqpP5P7inQCUbpg
Cc8WOy/d5VO46LjwQ3iUm2E6WY2nYR5unLTEX3ARriM01gPGvP4mFOrQh8HgyMDH/Dtn2wbJbVNC
uyL5Mvck9xxZ437NvuxN8izqPtfMKMOPRzFskVpjMoiviapp6lVEo0vdCaNMIbVSYCDp/rbOWfsv
8q3SSnKy4+zVXJyIOjV/royZtIXcmDn7Vzfb2FHK/WbBRunDGxUupvpXNfI++uh4YEBXUE2urrxN
0UsvJx6Xq9edu1oa9yHFUOJPbXLIIsBGTbx1RvsafvHeAeeT6oJyaJgTjY1BYROKMQ5hmQGG8Q+/
dD7/H0Wd7x62RO8jKYCm/DJds5fp5h7gCwRgbZBz/YAi5bQFJInFad9CJuSBC40Opvle3E8nkTsv
aKLmU5ibROCHMdsAhTtRYDG1AJ8pjhx0PdJWlp9XLmsoaGqmiwiuxPSzXoCkDnzO2o4qCT07ZzTK
fTSd3gkEgVTIsHrEUGR1suA2u9IuScXvfRJCRNe4dVQq715Wfdkd4Rm6dF5VGlx5+mj4H4WkzHRd
/Klgxg/hMQx5LNW/QbAxFz2KQuB90+buMT+swd0dY9eImZ2PQQWW9CZXMOuXD9SgmaGS6z/WkG6j
fif7Rg3Xao/Rn1KGE5qPFDf3DutAojU7a/OEr5kW1agZxI8PVw/96h09GDuFq9aJ6ZkJnGIKq2ko
rR3jc3clSs/SXZD9W9qjO5vc/doRNynMc5TR8cAcNqE0HtfN+e5tX5COJzNg1AMGAeaZSQAjdyat
jkkLElaL97qiEcO+2NXGzwXFuqLjFjPMr5ZKwZ/LEl775OOhdQMP2NtRK/Hs2JtL2OrvQR9Zk74p
ub73M5fuoZe6ZubO/HstoHlejEHTsFesOqVL6jWz79US7l8hb5SUqyJ1bwSAqVmuJQJ1MiQxazEm
B8N6mFpA1HtrMtsM2O5ZewI2BJXnTuUzyQuBRbn2hLoiTPf7gSOPl15uMMy4xPdJ1ehoVM8NmjLJ
+n1jvSBhtLNrpTXzaPLbbczpzQfJ+eu4J8JdfYkIQqgt5M53NmA8YKjtuQL25+YwXzczxvE6D1pi
wp/sgNojL4lJveLDI0N7zqqwbo4VjaRggTXWxcPosowQOlNPlpzt7c1Fre1utOAxTucSapmFSAuy
UNi/PKG/i8jMxVu9Y+iyEUMIDMP5W1LDFYxJg2ak5n3KXohaEZ+dx1PqS8otw9aDVsTwUYmTJQci
3bvAnh6kf2VFWSBzaXYCF/spOvdNY3yP+4AO28lj2cJcj1JCVkobFB13dRpFTwmQqXU2JPVctb+w
APjcQLQHUfoW7bruqYj2ZpyFPCue+Cvs757JdJFsvqOnrTa+DzdmRpVc/hbZLsPWw1B5scWX9nj5
w3ubozxNUEazqu/ONCv6zMOb6c5kPGF/Jvm+HVzZyXsXs6HWDQ10vAaVJTDuaJnYct3m5V2aIzFb
bz8SdAENIK6FUlWh4WCsAPX1r9IVDWKpVI/0l9KOGJeWsZ58KwnCL1JwYx8VSJE23/acM1V62DHD
UIP3bQw9mqI2nhZKIdapTif4ZZAiTlGfzm9bMW7ihUvdXS+iSRrZhh0agc+TYpyUNtG4AtujGL9N
tjBRIOsCFe9znkE1lshRODVhy6IMOdnz+uWQ+ykwVmz8umqt3V4LcCbB1bzhxaAqrkm1UmhPetSe
OdVecwzce4oIp68Mqqr9ASF7BwjU8u2GjuRi2+OkZW5woTFCjwQuwra9cA503/9jD0zN+QgIQWF+
ngc028N7MeVCoXcWQrAD5Hs59Y9Cye0Qwf5KIMwDArCJCgckhzS63kZYZ3ydc/vAoFKymNBgAvYn
TE3/UTzQhgEHXU6g6CkranvOAsbECdVfSihoY5yJImDCeaDbB/Ehe83H9PvAVi4+h42Wa73dhz4i
bK02f8xGS5TyEeP+IlM/7oPmKHiGF/cMioblK7wvElpz0RtYgcZrc35CmXPtoQmf96qHk0jB4JuA
Do4O4bYfq47rWL1A5m8FTdZenEahTKmahzOYTGxflsuVEMxW5Ji0WgPZDkkF6f3NUrtacaOztgai
KAY7cyihHfQt0LJfZt/RVdEosdOWtAtaSfxyudOCph+qiND4DJKkZEbuPshBCWEF/jGq9cMoXtqS
9b9AFhfVGsDUjEEGLIxsl/NnfREmgCWT4ltj3unQ+yEhvKyAaHLIoDIm9fxkqCwVrSzDxMYAwyrx
FHl2dmuJ6gS8Ln2uoOw5843QWYz+IaEjVSHsRHCencq+ZPIY1OqCLYae7/9y2Im5+RHt2zmTuXKa
51KXZJtlLt6ejxa3cLkUyqByGG7XznqkUwXnTPZXkqeWhu8zxZ9IXSbrJ0UsDQH+k9wHyoUb6Tgt
2ouo8pgNKJf8Q0UWsquz7851ewPzt9SqWMQ/L9ewEdWPd8zw/dSlo2jEC3Z6Rvoe8CjpDMovwKrT
GC1bue7Hhfvhwt0fxKeEdJF7m4wsnXTpUEWpDB56T2QBZPEaMLn/N30ax1j+h2iyJP6DUy2dMNrn
LT2DyL2pn0pwzHQM0TstgThagFAaWvuAbqTOFcR/e1lKSAiqLJGecf9lFcUpMTqC5SEcIacRoEZ5
z+Gjtwj7ay6Z0aH+ttLUxIZ31squ5JK/EWAprliwQuBc6fvMiAFkhzyN4gvI5UV1mIfOvNYBPyx3
6LdjqsDzg1OQ0C6/P6N0f4mMYB9r5MF1ZB1ftQF0EIdgc4Ckk2uWj8iN9R4kQxYxUcHYywdSqej6
IWH2PPbIklCmZ5LcOJ3MlEd7OXRJafiobFzt96MoiUmV0E/onxfl8uA5dOJiaB4R5I7C3nyOy1kJ
k7w78BBCOid8sN9ZC6RkUDxLNFy+sHCpsC8h++Qsec9EkrXA//FC25CbGSh484rJMv3DW7OEGinz
CG956IT6r+rbvX+Q6Zdr6XF8iEGo04cTSIqyovUqEzkIEHa+WXdBbKjZfFH2H87cx479JCK06IUw
sB+F/8Gq7FYxKbmEsuNGFSctNgw/dNjus1rQmBYh4RRY9wjPim7vxBMNA8ihem2CBGHt46ENIRDO
0jc1N3MmUFAnOsWT0l/EyUWMtXeXzQZdWSoAOT9epRk1IjLo8q1jq+EpSmW602055PwF+1yhan+G
e0db6VESjx4wl/NSThgKPAsAuRpsUKg/70lMvTL3V3wgjCZYuZ4nubS1EG+n+vOuKYgSF45ZKadM
FQ8w00O60jml4tsjXA83Ps+Ddv4z0EwE5tMsljQDSaIbbAgTNk39Aw9ftmMzvTY9PGSkkwWxf9SC
romJg0C95FxphcCiB1AOAtomyYhcGXk1qyIzUmRiDbmQTB5clUGHfLzopTz5EDm0VEadsc11+P7n
dF2Ej3T3cgXUGSK44zAbK711EGfMO10GqHxOZgf4wgdkPlSjasVFzcf6Qu2bUW81OHgnHcJrWWUa
F/YgZHCSyoKQPYuIUerVrIuYxdBa22SbzBVeU597xa8AVbpJIE2lTI+Fi2shx+WZw3xuXNZfBonI
MPZ0JNlMWjQRErQZrH5b22V+yXLBLCRyMJc5Q/M6n6Bcuvcp1bAYBeEhSkVQsnghyLAaU3qLhvFX
t6EOvfpGsKT9Oa/HXderTom5T0/8eeY1e6rb1g0xy0P10IsjG/x2XIgcx4afziCzhs3GgMP3/Xus
dXEteuTmLnSD+NUwT/cYJSVtmfgj9XzCKXKl/DIrEGlIywY214teLD+TMZnG8ijJRglXVCI38c6H
gf0KJPV+1Hv8mb4XhRjZr3zVnN3nVm99D71AKHWoe4LD1AJP0F3D2Wx/vIbqwV7UHBnKwM0PGfvp
hdmpmCcfn/cq/S2Iwg8ch946Yt6mRFkKldlnkDBNno+w95j5PYRzkPepwBR3A6hDBy7J0w4zXxoJ
+3d8Mzb3AZTe2Of65WWgYHFxVG5LBq5npVgMSZCzD/fr7v/ZvceuZX6vNBpW6LH5PnDskZhhlzd0
TYS8iTqn+1OK/uK/GPYcvvh+AEzWVCjFtZQdusZ/o9FKExJ29AL3ydJVT4ZyoLc45UiBJRQ1qyg5
c1OIRfHvT11T7oDj9elviLmr9sRoWb7PASpmKesDHqG5HSXdJH22xohh/ITWfd1a+EZGXoUWxAOI
gU2lhElyxGA7v/9rTfmyzXnz2BddX8fc7CizQifq/m9OuSis2DmcOCLx2SEQQ/Pr7hggUSM8nQ8m
qBqIaI8vp4FbUdUEzPnTpZ5Hx+l22SJVXdJXfnZnrZpZWrv+rYC1AyRLVm4DrOZ5Xz4PwGTIdHkM
yPPqPLDDIaE3ciYmDGndZiidUjLzxyOviN0fVJFVIy8FANDvabWo7loGvPpVHue2o1uvKCnIkvcW
I7gMJcWmnFBvCSNJrk7kSNtoG6rIYWyJCNcfMsKEYaUVk462lMsyk5G09+tRXMcBGRomqZMxPj9w
rPFcWa5VBc/oMWtiIFhiAz+cLRe0PrU7/1Egk/rK4Q3qxRrDfegBl96xabUFbGwItYRIXMu9uF7b
/fMwnIIqaxB5xDpml32u8t52fSJNahztDKjJA5/EOxRsAWAOTpxnbqfiTOCdV7DT68845eiwCB3e
LT0g0gsbGDKNkhGQbrDoSrjqV9GFouckcGynf1KafDO9qUMvVlAMlOdSBvJOJuU8srnhzQzY5e7j
Qux+iXIZlkMJaDByR56OO2hNl1GnnOa1AS0GIrw32I8NZoLmOve3VJZmS65RLjV/g3Xn6OP+O20H
pBVEueVyBWDiEsWbBvL6MpgOub572wOKd8aplVdrVh8Q0xUV1qmaBPccbQ6dnle/00an04HWiK43
rdqWO7z58uje7S/3mbo/bvEVS0Rc/Fq5IfttVSnoDk1SUpSSrbTE9FoDkwevL4L4yzQ8Rjua3nCl
8CecncjFvIX+SDv/1brGHL54vTeCIX5FsySW1SImJYMaPnU6CpCS1t0sjzbBtv/u6vouNMgu5QBy
YmB0rJfTWbOx/CKFblDeEOh9COi4/KsvjUCnMtiLLTtSDZEDYB5lw5OPcVj5+ntfDGuIW/ryxnYu
62wVX7Yqos3yC4Y2EiI9eZ3+FY1wx7AP0F85S6L36boeshTu7aa/ox78hgr0bWVBJFuPssXHQWoz
uXIGVlTLUxkcFWCwfPaH9NTu3+/25fdQzew+8E7l91VQaPfqPiCzGmfhv3WvVSMIrzBruDPnTiY+
1x8g1oRzeT/rAMKzpJ8uopmKA7tQr17XjDU+34ogcKehH2MN0VwnzWh7fhtbI+iuS7RwYxZ0la/3
9Qy8rymTXRaQOqvXt8P683XoDbeKf5vWxkJR4nUtczi4PlRBakmX4DLtQ+h7/SZunjYKzmW7tzqG
GWOYrf4z2MOULDPhwa147dMZEV2n/sq4WrXHvVsV+kY+OFKuiE8M6Se1q+O4UjlqYrC+ofM7VnJQ
CqY8d2LsDZtAYbdkfUVXl7MFlwSpu8a6OINOX6lrLB/9dCqRHOxo6vMmM09h98RK2APQEyxZtckw
BzbQoGRUYNv5vZM5jtmMEtRmcVq3bvBWngOKu/wYvxLKYeovdsvgrOuPj4DgrrbpzQ4nz4KAh14W
wmDdYq7Be4ILxBJE0emviRu18lrpl5jUGpxF0TbqYFqt5dQzOA0/KEV2aF3OYJdKsPn5yjegGrFg
BHumPe9Ce51ur0QpUfitmxsSn7fjRYMnbYb5qhnL/YNLo1OYRKlVUwwllO/ZJm8+D7Pwoe1bOjyX
2qUPV5EhtxYIgVQusZjG/Typsb8Es8brzWNJqN5LsMmrVQ9eH6MC1dI34IJhUYYcaxP9ukhZRH6X
nhAUMt+21nU16zagf0pqj+WPEce19ghjL0Op9LBOtuAEtornQAF4dB6f/huPrF4KyvpEVjCC2d5L
IBH65EKk9u32MgWB+LCjDVOVVsAEa13AausW8eHYETsP31b7a4FpaLecoa+AYUJgRkrwmNq6jHfQ
pS21AMvV8B2LqiMLYVXWz6skJY/zMLI5FfZVt8dQSUnuY9bbaC3/BU8w0pYlonecCJ0RBmzMZoR2
4Dabr88F0yK5mQ3JngI1ur57rfTfcdtJY8elUl9kIWjwwtnGEx4dQzJiUiq58xmKXCmpynQVySnG
jScGy3YyChhIiNIeDOdSHrvnjdz0SBSGR6EyXRM3kdzE6BEs/8lID+HZ4XZvu2e8U6tlYPW934UA
LB6dYqRxa3OvBNPHt6i1bFY6qjfRSGE6x1evwLIyF04IMxr55fr4oNkM12GEd+uOPAVpdvWzaiAI
9PQTtT8HLd43J2ec65dvpiOrV1Lf+ZB8MwOR1Ln3//WWacqK4IzchD5g5iCHTAEY980YF/MHWFxx
aYEcyNNPTxTROjgAozN392P4+Ls2Xna4ScTqyMjR93rTShN3qPY0FyGb+Na0utOkPRWclh8CsCoo
l+WcSFAROFnlgPfaIH1kUkVVM006O3KHUf4HlmtN0k92IO31epapCV1Oxls5w8g03wXsuOSBxapG
MnJSQLCpbN7O3aaI0uojUyrxwHhPVJzgkNCjqJH+GdFPcFOTr0/sbeTkRE/qAcCW8fR/tRAWwvIB
aWSPekDZzTydgRM2LZ6iilG2wd+WDGRCTsg6Bp9vPBATh6Z6lhQhwYpPEibu1x70IHU1LFxhnUdP
4eCofxikT1FBO/bpBCZG7e3PGvKbI6tRybOgI6mib8plza6eSh6Ps9oWxZPawYFmHQeEJ1TPkkvV
LUBIr4Mh+xDuC85Ep9lN8rjQtNkwK1IJ9Z2kN4stYB4xJVuK72EZTSWTaC6g/sKQcixTK9/HEmnV
idRm3qAQX4AXDcemDju8HFWuBCFXORddsf+JkuUojFfkaqvGod0OsKCMAQwheROfmdb7pjCGyDGC
IRMbjHRLGIqFqzTSwh3+FbMxpzFhZm8T3byvLswbSZB01ZZE0w0dTThywXNsIKQI1+hXkDJie2ss
RmW4zDTqMSfUKcUkYkR0W9F93tNvugvDbdzbPoBsKwihptiHDpHdn5aPTh8ub5dsV5kT5LDRYnB2
Ld40DyzsBx+Z9y2jdG0wka02IOqI59mugi5ZilMjxvdKx/YFdrHYSpCUjxgcZrI33YYWoUV+AOBh
HQjOftXtZ311pCqbI3lzwsVgcVdoyfZ5Cy2LSZMRVileBahnxfx8Ob73Yzg5BaJdns0X1OKuVxWg
U0LfRBQJHUzSS6GBdh561odWA7MUq4GpM3bm/BH+ZeU4xLavcMTTRh0u4OB1oI7TaBeF1vx7r4Uu
eTC9TD2unsEpxWjm05O6ACaWA86PZFznT5GfLQeEgDmu3mtZS+KwvnBeFWR9Jq3LFHYRnlsSrPoF
h8bTybZx/BWMuff8iarnKBJtAtJnJXov8CqVdzbyKVZ6y/XY+ZPmKo52tpBDP1kJa6vFjwWOpQPU
cDpC8jDNePu8QSNMtedE3Wcz75ZGFwp51N8xEC0BtYcgrzG/o57NeVaYVYTqlUIwTXPiRsih4HSr
4cvu/1rCQIUZAjgmwIazCG0nsygUYO8iiTZbi6C0mrwnij5Rxx7R06QNI136HWce1t8+fomg/pVp
mYngpsVTSrqeRC250wvh+iJuujbQGpadSVzEQ03F1lkvuAIzczPfKbcD+s7l3BpqqVzB98AJ5P2o
iwQ+ZZHHn9MAckakWL5a1s8FDZZlcJJwU/B5Cpl6FeEUNSDcHhcCZZu0coUF7HgNImOSyj2Yb1nT
UABn639LxlMgOmRhzr69mIU/HkSbEKwW+TYJ+u7LaHzXpqxfESEvG/d8sFcLfayiYSlJxgaKm7ii
s3K4T9WCbka5DwOATPcrtWpA+RUKQ3aNWIIu2gOaVvaVdFF8UQIveWCuduxJCSTyW2vdrmCClmey
NL+1AD1T7soUXGMYUNXPvlhuderxEK53b+JPuBr0by/NVrF1UskYU47CK4Ee6DWavg0dQIdrNgkc
yIMZp253C2f6hLLNhU0Zb2UCS2uk4RI6RbzYsFCKcmLgE7CJIBJwAvpZCphz7TTBB7pWRo+ZIepB
6ggxAwbS7V1ix5ED6sSiU21tG3aVyq1wl/toJpENi1iH+nxNjDPYazDhElLrccUsu4ZSccKB7WGk
TTW+z8JDh7/gKFL9+frJ6KP2JpKc3eckdqddqXz+IE9Qnh5Z1CBLgWjdyCM7Nrsd2h0Yn1SGqwP0
p6qbAecRZdD4g2fvKxZcRC+CeuQciMbS3BVRi61lamenE1Ddu1gLUMoQ/dMZq289B51y6GC36SOo
OMW+OY675j9nWXI0kitvs3hE3gRCkiTekodvlc33EiCL+WZi4fJqF6iZa+DfoRp1TFSu+XwsiRKU
9gP88+V1Wg8bqZRZdzaOKn0iH91apr0XioijuDT5V9ZkhMrU2ywTYn8kXSQ43zkfotY6jN+d2K1j
AtD171N5GuYSBag4f/UIe+YN2FiujGK7td3aFALgCA27+foZfQMVHsMmzq/lYknDRN7t9sSdXgvk
yu1TunIkbCoD/8OtEJQVK9sLy/AnLngd3mc7c+zyrt1tQaBNhuwbwYCQawJaS9mEOYuoRk4hgviD
u7dKJivUQOXQxLLyv6ogyL3J3/oEQBTEb5M3mEQNA2gA5b1v0EWqP5KDso8xEOtcwD+3A5kwB/ft
1tzYNH3G7l2PVXNTtVfuQgg0oDnmJqmOoAX9whfQl+TahIXRJ4odxk46RKNSxUvPf+zE1odmFkv0
sBOcKweL4GWhHMp8qAvaJqCz4RTPdlwGFpz/xQOvlgXRV0I8xtLx11ktNqCWML/EAIvMMxKOojVD
0B5OuoDe/W3+gFckxf0qK0rztlYWSSj62fvJLjF/vhJw5CN5wWu8N6dBKG8IqN4bXPBKU0TIKbfc
T7abPISVHLC2MWR+liN4/cnhjJP8a6SI7xssQjM5aTbEC5c6/ox8t1WTJPQLvksuiWXkrTBp6YbP
LrRQpUeaXTRGYaacsxIL/ZjBVjLnHExwnSTuK22UhmB2rERkrvnfifAJSBh8O0DDn3VaSGAiTe/C
OzEHxeTNR1Pa1BBycZ5B8KUSRQK9sOt5KclXbn5+TkJU/Ygk303La5N4DGb9oAQGUWoaZyS9f10y
FRMWcduZlBSMCkP0I7DVwJ9O/2QC02vp24psqFbkGRrqp0jihGUsZH0m5JQBAJ2S/MtbxPoNWuL5
xja0Sgp+S6+Bp3DTLODBpzjAIWF9/iISQ8B1YulMzIWNfWLA3mK2vYU8ZpY53YN21cQdGihU/zos
ilyoIvzXU9moUr4/EDXR4oJr4WFwTH8Di2nHN1jDPvJ2cVrCNAqzpe4tkzNQ96+Z3xjP27IofcRx
vrtCi7L/WoEc8qEiZ2hRStvCqG8BnoO74mzGIrPB8FTRtHle26OP8jRED2eYHkAex7QrkLc1GNcd
iq+h+2ZRpc8f737mdnuJyrMwpjD1RfNzYnLfzAXb7VqoFBH0rTy7DpfjtKk5c+ZOiiCFJRwtAI9M
0tgWSj2otclsMTR6XxaXOk/9QDM7wyOpSKB5yb5RZIZarrgats+zQOGbHNVStFrQwcJwrRrZCjP4
u2QglweSjWl7oUwvbLRhydVebFs9/W+Pzno8UYautU3F1fRX2aqaYcGnhK3UI5Z/M6me8w+uEpFV
/wXsJWG2AxmA0DkIyPn4+ZpAItTUPY6Vr8GT6BVNHYG/ADTZCxQ8mSaIfj28zkyq3x8JICzy6nfG
zsZdzmPPVNA9gH96ioQUBdvJblxI6N6pWCyYisiwMxTa5pM8M824vTV9TLtrFbZmdsjynTTtt7Ek
c2A3/vgVvFtDNz3kyC+wdTHa5mSWSGkqVIPmspVFDGjEzxNqNjjtmnXeCariXKHkxRzrPwyaWUi0
PH4IVeTgk+2uvHM4Wj31Jr9K85SoLM61UdEN/lUwegHC3oCxkhewfrgbMnMC+QBo6z6W7upkx7wk
qfWpTGVmb4WojHToZeh5E3D+Cqt6JVzThVKSVjYf03TP/nc/abb0Ow+p8FbpRNw/uE5mtCUh0460
f6ph7kLxYLmtqZYGW/EocpYWA93aMLuJYIjXGf3ubdahvuS3+r/v8Dhf315/V24UWr0sVHGGoIde
nak9N8lkMEzGOVM4jRhFR80ERIY+PNQN56y0xwcFmGf0qzm+VnvdsyAhBVDFr9Z9CyJhTWKwOFNN
szEEFMsyuh4lHs+QTrVTXDjR4hxrRNpUsQSjkBQcO7FvxYQwcFvPK9ibNTvJ46SwcgvHQXfXvA65
sF3Q4lMLqlhpih6ziRmik/ystGJcoRJpOMZYFCS+xS8cgymBNwFAuUvFkR2UX8YitcsIh0tA0yZC
wNR3kSeP5ftXxAZi+/cIkIaPEB2OydUF/ISPtZ9+poTU1qsNRhrGiS8rWap1cXjd/wfMabVFfeL4
iuMkJd8ZNmttHAZ5Wwzn7VlDY5A5kQ2Frl5pZYlrkEevbSaARrxqqiQ4N7UCsWEPR76Ph3M2nv0f
upmIdFWyTkNieRiCKWBY7CEAa383CKBcl8cCQGWruI9rtXAnWr2I+7OboRs5uoV62yiICmoU3nhn
XAkox60PeINa2REr6bEQ4kPmmhc6qH/YyiTL2B8/7Ly2y8gRobzrM5V6EV9qu2R0S9paiLfKQ6hI
JDLdTJqKavRXMDqH5ixqDq4TcoLSZ+ZIp4oBQ/GPfjT+M87xwg0XWrtgRKNTa3MC3QmdIHvyjqtM
OK+CcSPe06NLjyI0UhnJbMQHLm+eBPC6MJnfUGF9Ag4m582AtEYwATZzScdJN6OwzDYYUYzdfvma
E206ALZXrxhPhmF3pFgkSKZwim1uiFox4sagXQwUNjDVgPzZUpAmDv/XbiI7kebVubfBXE7Kchg3
v5lEpTO515Sc2q5PXAQ5If3ES8qCQksXJHUueFkssQ6nOFcbNk3H5LuiCB6apRZ9e32Hz3JzUkm6
0YN4z/4+EJF7/E+paCZcYPx/FLEjJU4SBj1+8LBfU0a3CQcz0GCmdmyOd6NQft7yisQbIt7+6hIV
YzJ3+lQ5WFz81xJp1gAgQZ8C4YUEkDZjn9djglO2KwNyKusUvB5N0WCiSmJ/av3clLOopeowDPEK
OkB+VsaUSgTJ73GXYhycxl3x01qdMmi48BLZ+mykNt9skinNGMXDqlZzvpsmPHk8kLMZXo/a42cd
U5KGaGEaco+f8lkM7aYuY0YWue9/JKbQcUTlKRX+V8CQFG1Al0I55AG6qPmweDdwCUMSBCqlxDFW
5xfF5zu/2EUn76kpxe5nyhcYdJTqv1DWop2hkhbc46heIN3thEMUCRd5GnrxcJ+QN5oc9+CQ5EQS
l3sDwBpHTsJoteWxuon9y8Zq8EVdVWJLks4sKKv5gMc2y9gKYrUeK1ZQbPhPeQiey9HIqSmeQtsL
vMgJiGUi7UObZyoa11jWnO+576WjruSFaHzUvJpov7Imnt4WVMRrq9BvKZDVoMNdWR5HonAf67vD
2LRfuuY+cFtOn7/UHSmboqACID/FmE8dwhFbhPY+0uB7jFAtBCN6XF/os3wqG00rlQLMCnwKjVI0
iwh1hOd7N+iEjTHzwDRvp3ktJClXTZF3ay8RK2r3EK7EUKOHKu7Ylbo3eszzgsMhVAnwIY6kQhuY
if0E12s8wf1qzBPJpQPo88yX0iG0kQJItawLbzVEffe5vTmliLv/Y0rkbx0clUoKeq57k17jUuv1
K7a6MO2dzLsdE19p9AUd7JsWwzC7bYFRs8Fq7l0zzFq/HQ0W62b196WonW0ybi1YPoZRasM10eEs
jB46PcukAvXYTtrOof1kZQHVcLm4dBzOPTEXaaPUEpwOan/3YLPaWyWjI1tOH3VZ0N5cQiasfad9
gC2WDRofSeCflKgOAwgShonoUmVOynRj9lVFyV08c7JGajwnuAuMXWnDJVdgWWDiwLhLXMj8QtDa
NO0CrfhIMnIl/D1tZN4C5hZ3RMSyj1N4y413bVcTS++wjOqneJ8y1OkDcpr1hZgDwIshA4jTeS5v
9gAOHH2im24NAITAVbBc3fUoSPomlrV+KvKjGaRQB6BjxNWcb0oUp9qcrWflkGxM/DtlXKbgKuo3
oZQapIW/mD82YCEZQx0qXNJrl/g3aquWMo2y4qcgVEe0MbEAXRDiPgDoMpLZiLGin8uMqSh8Iz0s
gYAqdcm4rlfjVxNmqE70NMst7djNj0z4FtopsHsu6GbvnExirp13iXDNSQD9fEgVGG3xgt5VO4R1
X4PLAV9VdNyvPxTHfvMxnhdRUNG+HodWAfwr6i+FyVrlQdJugZQCf5Pb00pg0B7wxtesYxDepp7g
8vnKe8dUowCTw5F1aof2b4TwaYZWYhty8oOFwDWjs7hPIxaGuzW5WL8dd5291nQmtr4DaqHnEq8B
9qedncNYXDu9CBcD5voaR7UfxG/5W6JdnalxuxKKhlCak+rIOg6CAU/lCCRkWxSVvGlsdiwg3le8
SlmbDrmWY5BHCcI/U4efca+3HrT0VjLbQSwBgMf2Fqdi298IoOVRnLJJ//FGP3uVRyDeGfOgdicl
ppHX+B9JX+bqIduYjeP60YipCyZl5yv9r5ykxgAoO2C5z2F67zjYql5ta6/nSmSO7Dp6ipBmjs3p
U0kgvodF4lrfXN/9YDA3NzQKpLtq3CH/Gc/Bm0UK/Fsw/hOx4qAeMpm84aia8746fqQ2rBrZtBqx
Th5CFO6tldmCvyV4KLTh0YfN3iqQSS3cCH1n5lvxNfe2c7DvJ2w1DbET391Cp6a+eFkGYXzRWyGy
EVUbLvwIWou2avMeOA+IljRnno0xnUKd3DoDU2m9LTiLiUbRRGQ65EHTYXZy1CSsROKuE4MQdK+M
YvNQTZHUpH5M7qDrl8WYkKh29ThZN3dY3S/A402SGfDjkQtY+cJEuWCFRp94Tfn3AmehiV2HFJFf
l4fnHj8bLDOZXfNz7von9/2eB7gXROsnsh3+QbNYmAnbTfjeEGTUqnRUt/J27rg1H7Tv4w4Luipp
tSsdTA0ZYJT13XkasOE0x52hWgh47GpqqDiH5PDMufxN2sNfr6EJAgFy10QkrCtzxtsu/1/90YF+
uwImw+RwPHfqVjXi6EEp2cVpi/F7d4hYLh2qpQWOegDoXOJWj+Ptw+ImZ9tKDY0dM358AciNIUhm
MZtRyrauWnZc3DL6s1ehpQA3R9avljVjTh5H387QGnZFaAyzprbogufW5+DQza9RNSzNyU1oQuID
/zO+nFtLZtqJ1eA73hW4vL6Fck30RNpiPCHd4GQ9kDyzvaZh1NvFgo3IOvQ+wKOLzkWzMcwpXV8X
0G7kRNl9YTmQ8M49E1NazytsQMpaAVQvQRRJUJru3jGLKZUb3DNlZikqhyia/EcWyWbwtmPND5BN
/6hei5FQhfIy6MbFlIv7kTrfWY4UVTFjmeFrZ0e6vL5cnVneHJKiKM1oLAJMnSktmtWbwrbnyqpZ
zkyUlLS4GmGt7W6NpM+fWROiK8SUlRtvzWs+9iyAeDoTjiMWYHzWow/fTla+BwBRKtztfy/mdpFA
PCKCJkIxoa84UrUZgHuc96oUp9xDPwAuGDSD+Lq/YnHvCxbvP6+OWi09CJ7EsqFG8lrIHxtqMNfc
JnbF8PuQyiBNnNH27Z2f5Dh3aOWgBSFYbcqCM7EyctUEyGgivMy4mLWBuKb1WipovlxFhyLPfWoB
ZiXWAqLpCgcSvdtgykNADyCUNvkIAkWEksIe4gVgfoEj3U9f3GluV5uAjZS3b6LBw21a4qQSQULE
55wyCqOR7IQSZiOzkRGpNZgrtSNYGSoyiOZT5Tt5j//OXWWRapGddHRZirQ5KmTnfKrIcoiyTqfj
qD4jV+sMOsp56Px5qdUv7QnwZwlNweSN2DdHPF8vH8goouqs4+0/I0Jx8+U0QKJlftmetDHWZ1cz
9knLKwR0ks6G/0M07UpOR+oJkN3Ox5els65162vsW2DHN0E4x8oHMyF1W3rv2aiO1frw5ynd+pqO
4+DiC3Jvu0+rTpd1D9A1YFHO99pmpd37Q811w1QwDL5FHQVmW0xEbV9Aj2Z4GsbzLgiuBKogkkut
iOck4VCPqyhs1KzuN/JMj6KrtZ+v41vifS8ygGl6kM7Bm1ytnip9qA0mC/dd/lzDqqfnTFS38jIn
Fd+eAtOCPXAyX6OkHHwZyaA9gLePgTOe+E5n7Aq/iNEzknphXTd7f6KEu6A3FfHmsKXDM9qOwvRA
w2lMWs7L70yQWVmuS+rs3r/qF4DvkuVLcqyZeivhAeY5fdnMQ7L1tlOGVjiWjxwhDJ8sM4kjwIz6
KsEZXM3XJnJ2dtdpZJzchva1FJ5x2NUo2CwSde+krwja9JWbjVmvfynLdYF931D3wX9J9mCrp1pa
Q7PsTt/cljrM9qV6CQXgvmqSy1ys09gzxUSlzlOuhZH0Ik00maIW4sQMp+wv5Bh+lZo2XqtSB6Iz
ss/45QCwBo02o488QfLkX5lkYcHUtaV7W5lHDNmmsEFVH6asT0i/ofIIs1tZYSLtK/MVddz+nz6N
SrOmaG67l4QLxToIPMDa79MgYOZIIRpPD8dY9bkQmodwr1IeftqnXAgGG0CenR+8z6iIoqA//xJp
R6A3ZTloXvjcfAQZXdpchGOeZ8aX78LxQyGL3i/xFvZI0xhctnGxT6Xqajd2LffmixifemoPRCNJ
dqJ5mKC9tNQyz8pSS7ZttTcfjIweGtk9Zl4z0QZl9lz6zQCV4Miwa4JMvIRjRnH/wvDlUsy69DgR
ciF3xFzfKcB266LCty+jyoWvP5YKlhvKce/gPou+3j6lJVhrSjlZd6Jz0opaqdCDNFKWXoVpa674
FsTSJ4jiub22dU+iSzFpu972H6w1YNnmPv93vSZkLBMFzsiIbrW8stVKw6Amq5WGyo3no2pnd2nf
TwLGQzlQTWKBkC3UiWIVsQeya/+4obKJv3fDY22dUvVMaiQSzl6xDq7rh136B8JJNHVaYz/o2Sdv
WkFkp5PFCwUJlLR+2MmPWpF/H94wQgLQENG8q+ZmGkd4gavKTqlOz2WoTSKllK56hxSmvEtK6YWP
q0eka2626mWmReitVB7uzgpqzBzLwt+lJFQwaT6DFAMLTVA7NJzclCkPeGPos+UgrGsS2tSEwzyW
bB7Q/3kIi54RvC2Hinst43VEXjFGxKiE6Wdiqjh1aDd/4ccF86yRNyoyberiWGm9g7Es+l1WlzNp
uQwJttVdKxM5pb7F4xbnjitSeo4cLmR2heX3RcXTN77UAqjL+Jsk0mPtQj/Dt4j3sjraRrJr1NOs
OUie1WFNcqav1dk8yl+GNCOrj94yKS4ALRB1Vwja41jPKAomINgwK0xWLKKZQYX+XMzjS7bKFLjd
pd0b6nF0+4pJmXCqEpSiYt8IU49L9P314wecpiQcBKpsRkmuLFh5y56VtW4Oq6rwdtmBPKWUP7BG
6KD3/e/ehg6EasVUeql03i6RTVua2YQdMnIzLgEC0gHB0+HQJTFrny4XhLO/+i7TA4Si5l326aqy
B76W9VE9m3zqC3DcPpczSCTK1v6S39jmo4P2KnpcQL5WHvMbi9m6nrgrM3Tlrlpd3uGOZlioXb/z
mUSVOPxiINvsViDYCg++m8+hRFESG3Isy9vYmAl08nkbLMr1BO1+vUy+Y/PXV8kLAuw/1HBLoqmc
XPrs/ts2gY46hjwiZwbMQNsiIqpAgOyjJsypJMfkwF2IK4rJfypXLpYR8sWgOS2nAskJrSO0UXHc
pjEEIlmVpJIpEF/Ya3Vr+V3qpMWcK8zjLSYbEZsyQiq9iPg9NqfvTKnINA8uTq7NKx+DR8AHAP1z
1A0n1ElYUBF+SeKj0RuB/Lm7YtRZ05RAORee/a9MhIOcVVHmS6dDvT6dD0wysZBs1O8Smn0ejg+q
O/7Sz9lD76UMhZjI3R+d4LOaNcEpn4wAerVp032FEnr1sLYL8+FkX0Hl5EWjdHZSXCY6YZyD6QkH
WAldP64uPBburjE2RenOQHycf9z2UuvjA36CWFVw40H1lVmL9tbdSQtiqttNZdo7qfV6uM0rQYol
dQ7osA1PfVBpMscDvDAgR9IgEkW0eS939GaB3IqYXq7q2YclucguG4+ZtTHyz6a6LGz5GDGDuoKO
2fE0lOn0lsXv0TCfsX6iRdg8FtytcwFRGq9WSVjTXjTkeOg8IKc0kJwQLzQcrCdDkEQsklTc3hQ9
I+2RJTMiD8An4Znq4V88nfcZvfe/mS84bG31yWZs3yT6q00lqx+U5tXKhYq7eqWU612uV3Px+itk
ly5/SDBpZZ9ft3mnTjZZkIDFxvb18RsqMH/D5Shr6VWkrbEsf/f/8zsUZ8uFd1FrEfSIIw/1SDmH
hSd69GA+yet/briirSlJXPoGfwg2nSMaL0VQFi9M9UZyVIyLruMExZ08uSmDRfk7ygvvuvxhHtqd
IOKfTMcIhDEvS5ziIm/HBMW8v+sruRZOEal0tmjxxWOuokYamRWFEs1VWUruiKKudsz6vMaijKna
f/12UothljkpUSdQGrh+91J4NVRYkyAUSjo3aW/34xL668uoLR2xYwW2fg14lQOYOf6/ovogR0+a
Cd3evizJYtVHPEMXUZsKDyamPHno3djrEwNJhtl+E0HZ021dQNGkuckb2pcIHvcjPXunY04Hufw4
A7SJiJ3GlkaWsmZuyOW5trtZywBqIKl4ZkAooyXpDMD8hP4NWyfSMxd6q351j/+AR84uRGiXkU10
c22qQb3SMWOW9KYr5gx6O9B5Z3UkAQoSlAAd5Eg5BTSTkJXGgsS86c3QrMgShHZXFC6/bJTXXaRS
8MKxG3cbaCxxuPDRGbzY+58etmp1gDLjEdqb22heTNe7UIsdvisC3arxLNhwuMybFjo9VUAcPeG4
l5ECU/9g6GNLP1GmcyhWmz9S1DsyKVzkhJVm0kiFopivUp/NZyk5aCAqgKrCRZNh5ghtUBUIOgGa
CeWKSYW2CescIeFuJn8uxz2C0OHx6FLsMBR5cE7/2PxsWFi7DYc6DVTuo/XPX5IvV3jVmHxqA6qZ
bHze4DD07crBpf2bi5coZ5E+yvfl9QtOJA4jfelfFSpQCxoMsLyKBB1oAlo4Rk6bOti9ftHQuDUs
JHlhVZFYgh/RLpZiZJ/LOkUtBLs4HYeOGAcgL2ffNINr7kSn0CLB81kV6ZgEQLrkGXP7RJk1jVDn
JzacBgCMLlNZpDIo0yHCOMLbQDgEXE8RoJ9hNmAqe/W+xtkpTku0bHOon4hIQL1/D9Cd0fkj6bSP
okUzDDxQeE/yCoA9PwKiPiijohkSTJOt/v52Ib+JfCzCBpHiBG0zYgDHRpFOBdKZfMk2yThEmLb6
9XEsn8epdvvQ3AtI7hslmhAcpZaQoqNzreuWFjOgCNbFsgacfZ1C6Hgy0icEU2c9LQSEBTRl8Lta
9d6zY/tjRpDssxU25lwAa2c9EqR2L62VgCYWWCF3uFLIpjoP1o/5d5RdKbyiw+UUky8bBDrZDrSW
J4u1V4NI1adrdO5QClyewRjHelDCLSWsSBhwaeFFOMnjaWWOduhYMgFlf0boyOs8YQikRsmZ3PQL
WzHl/Wli9vRJoAcFejMKSeuvw6t9pbT2U7IfIqV2oMtoRtBut4UlxUmb+rB0SW4Fp8E6Idm7vXke
W9fvcXQGHFyaJDT8kEiqD4bwiLzhCo0FBkvgPCYIbXXaFzmiFGSXwHyT5C5+0kOt8DlDgrSUMGgX
vXS8hah/0xpY9s3YN/JDWFL1Th9BduDLBx/QRzOe+EJ0ILMSz5/igzfspqzx4ph9Wy1nva9CQpCi
p1v8iOqkYr93UiSoQtxPm+C0JNGfPUkG54uotdwXJ+w462SIXwaZFJ8AY6/od3JkFSrGdfK8APbI
B97qityxv+viLJAGm/gszmSKLjZcw/nmkQDOwOoniFmIq7lYqUhRUaTaz5PdOSZnpqjpMQe6dxFb
TuKXpB+X4ZgxGrqmpx01d9dOmV283LOnlVgrSbF9hxg/Y8yCe8trKjpNgAeIoa3IRiTuzQgYCr0u
1bdMPls83kYw5XJSFDv+Ab12Iy978hJHP4Ry6k5ex3/MWc2e/bhTTEekXtWWRqQFkxhvf0+XSwIM
+IwwWJKfbyUM2k+vIFdBoCubugjEFqDjRJgrZNq9q611Sqaen/dABlC6kh1So2He5RhbFOyviUAl
dcuD9iNLLGhgBOLuryluYVN2hfKkG+rPvzbACXSfr4RfTNgd1Jto+E+9IoLVRgyyErDQ+qcNatt6
ZmYKYOgBCgKO6Hje7Ef/fsbJq31IBnYHSawyePX9kA0+eBXpMQa9pRqBEIZLZVDB0M9f2SxcO7b3
bDBN5/l/AQN/SMnk5WmKWa4ll2BlBUJnYLxK+IIQK4uLfp1aBojhKayMGMco8mDAsPZC2aQCB8Iz
iPAuosF7fpJCgzKVZZ+SlcActgCayJ2zokrURwMFaOtvQx6/K/iXH1lzU1JtAQ3pwGjr3vs1lSKz
PId0QUUegPHMhk6plCXnwjU2wX5KarIRNoLuat2TsarlED9eGly0S2JYqcHUaX2TAIwcS0a5NLEM
8UaMBOG4AQy4VlSrNfvVYkNmtrd9/+wTj02uVkbaSXxKHhy9NPOgigoPTHvUkEK3mCCkcaZqOvcu
nX3Bg3mPSVNv6P8WK4rsiOydn2wA9eScyEQDYAnTufPlSx/2Ay6qNK7bWYZvGOyqgvrWONe+/odb
LsSeqmS1Ddv7LJESgrd+x2+sRWiixafCFC5luxKS9qhsvsKg8VShIqY/RocwJqXyO9q3j3Y6E0XH
mQcVVApDydcxRZg+M8Btq6FB9WBnrm5X3ematPwmeqBC1d7cLV3tXkfE5+8BNHQHA0GxvvXnGgMh
GgzQLufLBmEHjILivDLzjIZUcVNiC447yzg9wUjb5zEVGX66CjMcPbROyDJCF1TPgW7VlyJtL9XU
dQW2SjuHUeXI1Xao0damvCqPzLSSMP6fpvFkC2S1Xz/gjFIb2lElLZv02hqR1K/W8xaJUM0GuvTg
vv/nFuczG62q7RAPWqm+Yfs8h1myLdf7UfxM9YjwjkC/aqfp2Hc+PNSNSMDTWdYcT+aDVptf8wmK
GAEbGyUw3lBsdftIyrxlMazMNpw/bwBqif7oZBtCVa8FqGplq/YEyUYFusN8xzr1hE4RRy1AT/bW
jEqPaK8VWEvFS0kkj6maMaltzF6bafReX4s0dTmksxh0c40VKfQ7M7LiHG78z/Bke7dDlc4dkDoF
vv3b0Nuh/jmXMsJmXyk2J0ueS30iqcMbQ0IQSDGTbKGC6KmSyLtQOMhdJ56HSQRzdWWD7rRnod4r
OkwyqIgDnihXKE0wZymbgR2nOkjo9yMfOtCLRLtyMuFxB9dsSptNhGXe54rR86euhZji9yDDtAdg
YJ6bMGbZWbQ8qNMAmN0VKiYKjvZo8H6F/GyKeW2lf14rci/vdrI/4/IHvgXQ6y28+6LLvRySmxkS
jo3Ach26iO46sk1+aPfb2GDxOdAgRHqr0f3UPval6VE11BaNdZyvRiCPJgjr+/HOL7qROaH97pxC
a4scuCA24uGsHO5EH3OXqgcdTFvl/RBcckOvTS3+8PnQF0m7+D2uvllUNBdX9PnTwH9ZID8jkPg6
xw7p8V066wnIDDCoCe4Shj/c3RkuQwD0Z/6OB61JXF7cIESsMTXxAYL/zbHzFW6pYO/5XeMoU/IH
nKvxho3J+0Q7PYi2h8DucFq8fyqeRdx0S40PRuWE9qNKu2OfHELAE30jbvyyYhmLgYBxUm2v/s2K
Q6PPH0olJpQasSIsande+BlNE+d5TOg+kBxO22gp3T6dY5gwJt9QvvaFVL7n4MUwXqJqq9bTFPCm
Iwjvy1RcKyNNoB9B0AFLGdstzeKrMPQMFIqwHTueFyHzupPv1VBZhCQ8HOJLOwXIqVI5AxgZy+fv
R1KHcL5GSKkWv8XBiJZIJ4vKA0Cq2R2884L28DduR86R1BKKJUlSYR1vJGxL6lCEtsL1ZT3rE88q
hQfAAz9jOmzd5CaTB1QXkmbWwvyhB1rwE5jEUtUDnT77yRmKBmsJzC1Dc6tgZe2rdRe0+LojFsjL
uL92PdWAmh3KWO6Y1TFtkG+gtqDcl6jMd29fLsmOovFz4yPTZgPwGIvFtWdUqFYGyzVLrui81s6Y
s5HeZCFM8W3PVNfHd61Te06IHL/C6ZQDVU4NdDaVAXJrfRYw8TjjMRRKe1/plgapbNDE7jlwJl4w
c8QUmW1xsD0i3/quoISdTJ1EIEsnt16fD0591DYzrD7jwbBN5zlJjRb3ChhIfL0dP06RzBUt2ZLZ
VT28QlfcEpuB2ZO/Q4Ko2UsPx5HmptiRKAxrqHg00TVLR/itZeaTcUOTLRVUoGXiksfQ1twMhZIQ
W1tF3/qwz31y3a7UEdI/9R5GHyCcyhyCM/IjDNwNDlOJfa4CoDEzbi8tob7drLqs8Cs7cnqMxXI7
DOzkij1Wh8riq2VTxqJrKKQzNDNyP0vpWtPHOE9e7s0B48QhyWpmP8ejHJQjFuhEjwlWC6/BKr35
c8gSx4PiwhxvfOWL8lBttwU0vTqQk8VHEDCc/DrrgX4otL2sDnosFKBYvhqpVTg/rAON2wkyGNnf
lwpLbGDjEXtPtS9JJq5pPluPxpdvbL48/XGpWDJ8ZwM5yBB1mKz6xtYDYrkHDbYpO5KqSa4otfdL
lWoaB6t2J2IXroXhkkXfKmnIvNBBJzOq5Q442E/KMgSNp9nWa2JoYQuC41f8Ug0MLXCTYYysHrIp
ukmQwdHkJ8mFByu/6aDY9RUKfFhDrwTLiqbIRU4uZVao0fwqNOaoff4PRpkNBOj4CAgO0E1BjYIu
6+d9yc+m6OGgWmhh+qS+1vlFp2x4AjqDGbwibZGblbak0wa/7cLdKaTSJfSLdvL63rxikTtHbbPE
4oFyh8YqtW8SKHn3NOZUylVvy2a7YVjLfc5eLDLHBeThUH8po5gBnvXRt8ZhpcxrLPQcAvn9CWMt
KqNOYRE8K4OeYW9gOcytsZsfdwF/ZeVbExIjEkdiz0DCAaOzP3UkXQZF7MCq+UY4P4+zBAALMfU1
i3EmDTTpDZj0qNM8SOZzU0R3p2AB307j6AA1rFqBsuFK/GHUftjy2U5eUmY1HKPIC8d/TQ40gGdT
2/3t1pfwj0wwRUPtaaERz2YT1ubN/rnqjskWSbKmk6NYip1h86y8oTSybtZQ0FL5gZms70Pe1GJ3
lM28dgP8WqajnIMJOoSVqJFdDbQCpNQ9Q2ctaUjhwxLAz4jyI1xJAI4fd+hWOicalDxoRI6p0y54
hW0S1Q6PgvL0VzOAGjAsYNC4ExiUKKPfZCdxqLccYxqIZaY4XrF4ZZ53AR0UG/DTdCFu9vUhtXYy
WYzzHWYn6vyUdHpowJ8BYbMGMiw24Rq+0bMFHRxuHPb/6s/Imdw8fsv5pcj+vNP+0gJXJsqJBRnH
xeasdZHO5ivsDYM7bUcuQxz5b2JE960Se2ws3mjq0h6nuOtL/LE74K7ZtxBXO1a2cxAjZRU6myEN
1rRzT+pV9GEwd+IKWPujQUsjE+FNtqv3zq1hAIoGna18K1wRzr+wX/DEBakG723EvXZx9e9Fca1T
mDWa3pTF2vhxPd08F7tfW8t4okxX4oqP3hJnQWKz+Igz5tnnUR5UorIrZwvf6T6dJwHtQ8Lk6JV9
wUYGhPauajildxHag/mUpqrNaygdpkpZYW8LbMWk9ZmsTr7yfa9FMb83OEbAcoqjpOw8i6k4gX7p
rzfSL1rz9CfmA7/lbj65LEkekP+qcaDTZRmkKUF183Qj7lwYff7/vRsmYgDeZSJJipGTJJmomKI6
qXUC1lge2NV9TZ1nC/0eJ76MyS+UwNcQN2/UsAS+tjxnKCMBYJP/O29z44WYsvlSq0u1DJvZ+i+B
CNl4hoUALoJsipuApFwxXXwtAf20FMRNJ7kGWM6Jr3RsuSZ1uYzaC9UsowmeEgUBvsvmLzhYpWMk
irbpmw644Q7KPhKPTfbmjHmwQVWjcQdaryJwDu5qlVBRaF0J8/M1WFMdsBtT38bf2bPg5fcnDt3x
9jKcOgZB7gkoIqItLB3r/u7eKM7HDR+/DzmGokVXnz9396vQqIh8GkFbhNmV2N3eTynAxQS128yt
teuRwLRF8ZALmz70CgU16DVjxhv//fsyJ1r7yjBE/SFq2VNMwOUxyQogpKhle8JbtVI6ycl2yPzw
jRPAiXqIyx69B9GdKcJaiO0Zt+Pn5IMtYSEFGR3DoGv4WkRPq9XV+QzUH1t0uO4wVHQZkXhAKU58
h9J8bqPtYljVwxd4JNYUsWybK6BGfwTCi8p011RTNFfwmVLSv+puw56S8n1mbTYovb8fKL0JaWrz
c8jdTRuw72oHW9RYrGwrHJaySSSkA1daNnLin1KgN92yQ5C/By1MXrOPlhDWCkP16KEnJWuCtwwr
BCJ1b4MUCqYsjTdC5sXGWaW7GgIbUih7kqsiF9UjpxtM/wc86dVxO3HnC4zaXZ29mSQo9j3X3gRs
zikaMWCIXASTyjMoyeGHy5lm7ILxh1fpNk4Wrb5mY17+wcGIVGV5erqktX++kKWS3VBEizHM/9in
y4+8Xk7a/Q+dFfDsuAInEMMjtpg3RNuJiy0USdUNqzSPhCMDYNntiPQekh9CuBYg8Gc+khO2N5LB
j2ZjONpun7j5h74olf8h6QKnW43FN4lr8DbO3LKMPtcvl9h5MsDHsooMRgLcY+EWxbtyhC/1CuUE
sJHBVaWQP6fFsZa4PKaAQi4VJ+TpURqsws/V14tc90m3CQRQWZLJ0EJPAX0P1qguGkSVmwcqJ8AQ
EAdFCCa81ao+DXN9SxC8rcs7Y8uTRfyqoKKY3EjMqIPrjdumHuf4xZw29EummWrZeTCCjg7SySLG
Qf2opj5xvO0zjJlVAJ677KXbr69x8uIEnD5FrmuPgFlflgzjSWzGZr19evyzyoLlVkI4daLjJ9Fg
xuCyEApK39uphna4ouJ468OtXMCSsVusGhxdwGm5mGqRXt0eha0N8bG9nHrrVC9mtVAmYqoZchku
5Vkt8h18FU3kOnK/zp0CgZnF4VexNN2i9Pev+q6ZNZ8maA0KKnY9zV4aemhjdELcyvd9NlwbXoun
o+cXaF8X7CLpZskoTfMaqTWWlnWftOJJefaGMsefK2jBLPw4onUd5AR/RsLpcEZEj8iF0vXbEAKD
joIGU12inIyJuOmlkvYUBoFr0wNX2lQRYyptThz3frIztRBZzDYqjcAKusEXgGodKzy8HWRAueGb
UPdWrSfLtBkA6z0mubXnnTXhizonvflWdBzZkBnLVUxxKBg/hG31vzp8wp9USedFPeNYXaXCCqzc
1S+K6U5hl7nrU4OgJqWfHO1z0Qp988TAF9n31xUMM+yi6pX/S8UHTdb2ycc/XisTam//RElP9Th7
2KRk9cR6iQlUZh5KLgCi0S9MXsklh+HuOMOXMYICR7wdqZ1ZdO0axj00FYPUMHOJHQjgMlKXb1aE
t1/5s+eMuWKw9iYCQ2xIv5gKDY3dhpcWtqgQzkuq7E+eaDRMWqoRc6BsvF3LT7CiE9aCk6Z6O5lW
nlyNIVyd431Ndajqr2IrBTuod20jkqI/0mnjSxx63UIp3nVhYetq+J94LjtjWUpRclF63bbOanco
KCr4iCkWt4WUONRPpKoaAqR+58AGzkhv2zxc2sd0se16fyajfdOSHaBNEKwGmJ3l+KExgFFdAa/s
hJ81Q9w1LLIbqd+t2y7HYoEzi96i8LLcDUlNJZOqsGwxrRdoLwnLtnEoj+HEzF1Kdt/2D6Zv131l
CVwFBVNaoSy974QYuEBJqAXjiLRH1kvjtkP/kjGR/a5MGYCpHHcHz2r1nr7l4EEwkKKSSyoA0HWM
8ZBMBt6mMG/GRiqmDmgufNL+OBgIKFeX2V+PG4MezuuLpuvQKkEkQIcHuWCkJB9mfN2mytxqLpAc
bTkzLJef40bkDn+krakmBAshgMuhK+dooJYCek+wKu7NqmX4X0IB5C1C65fHKT5WV9gg5+8NyaNk
krgvUEcikFnUJMiHTwOxpCdkzTHpUPGVQMhe0eMBXAwUjU4Odiws4ehz8x7Gok6wXhCQ660fcWYr
UkwoJmPXNRnjNLQANjXQ3CaOQUiJFA2bFT0IVv+/glIsFLqCIDiTjzFnykUmdyK7C7U43fO9BjXY
d4lSuOzMLCjL0X/g9n+YmDiIujpZkq4MTO14bbSm3TJvQRVSDUHGMsaZY9vFjQpritIgZ3QtJB4m
G2XT73Y5ib/PUX6OhtJIO/sRxw8WwGHjWcu5uh0WjUCmbdXRlqS8p2+A6zmr67Fkk1GfZLjAZpPu
9QbaspQ8zenTSk4tckPh4ol1SD+dpnULkAGy/Ya6eJZiaUyK7obf+WrrwUjkXBbFX40gbUo4g/4h
ga+IUhUNosDNWFCZSvLiPTKd7BGFOEa7aCAR3CAVqwHCw5NfT8M460ejCPXl9ZqpMA+m3kb/SyDX
PpZnHMV3vPYfEE1PZ9i50l7VRdZq8ijrGtikVxl39fXnIFgHJw+ZjZrQXXSpbHtZwESrwVYpuZvN
UKFCLaZ3Dd4+sJ6+IRgTFGiaT0TRBixrkLykY+qx2z6d81tUaVKOFmhpM5uRcC1hUXvzRCHgx30+
2Gi/CE+ulkogBzTvTl8WOhBtFp6yF6EDfS9f7q0SgTOvDGoAdi5qkQSG4ngVv9Ckp8d0+z9h5QWI
Tvv/kfoGXabfDj4N/ZmCJZ3rh6oNwykym/5KYTNl/bhxB7SQCiekK9/QVgRoCNd8U8w6skNsFu9m
MnatHXIqXrP8Gq+mC6LX5moH9IqbbPIJsGD+Jc+m3YtFPm0fBw61DVun+bdvd7ejU03Lodhj1Uzs
hNy73PkU5+y+FyD4UWdJLVdZGwdOR76gdJcHWaGGKm2aZLVjREBPyyRp/WCyC29n63YJaitDICsy
agif8YyiEXQ4xmKWnF8v5dgB5YAqs9TJCZLf5js6zjlJY/LJIxQM2+KOwgi8q7uxf7HT9GFUx+yo
RJTeagRMoYhS+vwQe4zA3YI9M2Z4QmpMJAJfdCYaImBeopx4KqAyi1wMENvwkuk8ZErlNc6QBwSa
LZeRbM3LPyPjna+ZHEROGBbkkuvmu02ISV0q5L6gy9Yl/Y2uw4QV12D3GL5pSNWVuGQhMXnLFKjz
lrIkQShMJdL8WszaoOR/TjsVHI7NGZU/55zbMVyz9K4OQ2cAmhkqp4b7fMH8KxTHzljN6B4rifhY
dKgoaJ9vt88iHf2RKJR+kul9IH91+wLTLkns8s9egao2Wv4C3MJEZJnr87wBeqwTuiypETlnonwH
pxjHsqvaHxYWOFFRXCM5hKRBJWP7X1FQlQjE5tojNSQW9NvdZ3m0HZ4mQ0MYqW4l0bhNtZB2KxKk
bFWOisYMvcwXEsJf3IU8zOeYbfEJj64OJDs8M248R01vxGVa21B2PejGgaRbOP9A/b4bS8e9AWvI
rnIti4yQRMLRZmloL9IbAJIvnGQmmft1fPAVP8hwJ3X4ppKoFe1e9ef2GuAALjIkV9085mawzPoM
Wqez9R2KVrzOrbSiFS317mn4aJBkJVxidQ5KhYZTJd5wCH5G0xuawXHiwRZteFlFrKjMLpX/ERy4
dMLHiI/KH2dI9xU+O81BW29SatBJc9tBJ7/EHRmZWD1EGqpuKG814ftED8zd5BgV+wvquX0wVRM4
7jU/pYUbJxUTj03mopDbaMAEbEMSzymAgtPzV4tJVuKBWknmNAJ8S+FPu+Fj4XtAmzkS9DROIVBJ
ePkFDXzTkCjFrYQzBPWp263YyLwdn0lfc6VfO2/T5Fki//kntcuZGRGESbrq/TUKPaBzhtXWFxbM
hVz41hiWamIF5G8RIH4XIBgtVnWNKMr36PfpNR3NORY5jM05/4eXgi34df/7TKosjbC0fzYSRqGy
AhWDn1Jvz/4iaAq0KfRqfXKkaNzFMpmtNSsqXamYjTgJtAiX3gXmEUZZbSR6AmX4nyfA9/eCArMk
VMVg5tihC+m1rYPX4FyO3lu6Dk7mbmqSRSbKwFL4nriYVB+tAmj7DrtVir0Y9HSdgo/6j91nqtuh
ux0eNHMEIkUh2+XgI/dw6ZGLCOxNkAFcVzMVxatZbqJUhI7HUHVuI8lXMQEkhCiZwgG2hZhKLniJ
VbCn+WT37j+6VSNd+dNlKHL4zh1Su/9s1U2j4KWayPyu80E56PB9EcpAk0A+3UxhajwHwA+DFXe/
Kc+3Ehvre//RbUZjghfd7/E5vZKNrWU+UNBp8QH0GJE431e4RM6DtG67RaIqzrB7mEOSxrzV4p6b
Mv5hALvaISUBPnil19TeOCgnlZZSqmpqm5kQoFAf8dW8NqWCdhzX5CPLVOHamD4vWlN/bFIOS1DC
A/bOavhSbQ7/yJ4nrJ//qS8wfHO365B+arltYwGXFDgUBBR5w0Y8AE59qDCGkzQb5K9Nc6iS4LQM
a26Hv4rcaWdj9vfR3APxrYlFEYmHEahWYcT8/XUKfeYJeX0L5rZbx0gtzGQBgz2UgrvApu5PDOn2
5Cs+JWYP+R/D3MD0qKOVltKewTJYxAjFm9b+9dhi3gcDV0x2prtqn0Y/jLQX/iy64q8oE8KqVcBx
UIH6ybb/m6zjBFAtUTkMVMrsF81xQpu0dknSuqwcN8D2hEmmpiCg85mL0Hb6tW52PveTBf/lQWRY
2pPYEEOA+J1ixMJDqyP2nUeO2/8w8sTNSB99OEixVe0k7EvWIR5QvVesjiAhJMTQdD/9iVeWZ/Fh
v0FjKriL+A7W4buCVk6ScOZT9C38oxZh4yncN3yn9qkIUaeYbvWV7i8EEkNTEbeJtMS5JlRs7gQu
kKcqR8VYlE38FbdYi+S4r6BeRNzs67Byw/96BOT8rgWULoxHfDdYh3B7ItnA5uck/xYrL24Z/aAf
ghzTCp9CJExmxeX36UcqDUOSaBYEWEZOcfqr7rxIkmyCncaa4V5rdEF7SQgQZnKaLcEKP+8DdCuZ
VbF5FXowCuG3oByyuSBoIs+kUBjcZ37IgaSI9dn9ldYgzEoHBkjVa/ijHc9sCHciBi1UWf85/N2l
NiMO7thx7mQedlBt0IPZkjGJA5E1QGAPScMJ9lTPqmZ6Xi1KliYE1KiW6CxdS8xHddHnLKjwXliW
8JZMFiIMdwPyI6/UPB1xvpyNGmka/gSpdJqMMv7NJEfDGKPEcvdD0WZgJHqmnB//z4ci+rkLq5D+
vIePpgKRWsYn/8YYe3QJsYlfR3azTevJq/ymld/XHqYBi5g1EmktOcoROBohfq0EdXh+BdF0Q9iy
sosDsyl11L8C57XpHv2Qo5esO5ROREkB17dHm9xO5yp1/yJrZZdPWyURnDdHC8T3hy7U8MefVqmc
OAEcDoSQNMS43bGEfnFpOcBJFYhzvEJJ4KjZ750qNbe2lDoPcL4fZhGDNDCviERUpidxTAgyU0Bu
lQE3UrhB5ypsiXTSRIUXj7u+GGE++VttOqH/w0VKoJDELyHb6qt2CdMv9V1mkOEquoBIIhxImn5O
tFnqrvJr6v6FINWbxKrw+wrjPG1CqJY+p3lPhc+Us/4YueI308tHI8DCPa18ZMpr9LpeosXhkD37
rl3bUSC6bzewR9aU3G15d1Z7YQjDEq9si1bYEVyWYttfYUnecGTHEetP3Hp3s6C/GeEa94pnlD6a
myJ2yN5AOT6xIGIRlSOSa7jqjpak1anjKDVKKfWYLgkVRCeY20XHA4+eNFfK+xK9/ICjaw+uD+PF
vUr7eQ30bJ2K+E/K/qjiW6Xhh0+UiXHPQJrywFufVTNrAkAABVj3Kue7Wiw/34rHzuHwpQ3TL9Nq
cUqIblFHEsCiy7SSiRy+FMN960d0iPNB4NfoJGO0q8YsuKmdb/1fYj3tX8N0AJ4JwTDMXaCKdCU+
d4Iqd8PlakheL0SNDFs158xfK077RMxRpS//TZucl7vfJbqOhNXBekQHN3ifYD082dNowTsHE+5C
WddRVcDsyCl4xOT0pZxAjKHCWZIxQTi0x+PB5mq1eC73a0xpvX2ikMK93RucEKlm5MPSvhM7TYNO
ydxKJD91l9O21VyKamHS+MfRVGrNloam33zSUdrGmIbfbvr/ugKQiQu2JqjAs7k2Y8TAp7dCOZxf
CfPRixjOPpx7k3GLHZ9/XaZ0W48r/VliNoVohvu5pYlKW52Z0a+iaOL85D1DeJsff1Ct8Hndumac
c/0s6RWRA3YRLIwysn3g1Mbz64cLgZK6PkOGLCoGd+55m666c4AGeN62+03LosrnyLyAIfYvRHdb
2qBp+Bt1lZqML+51vOW24UOUf5OQCq5xpShBsK62PbKxStwvMSul3CaETVgneewl6em1bu0HgMSQ
IsDP0kwnGGSkvdZlTJrlQPJ6K9awgRClCUyeEQwkLp33RQF3YPIJ4H76dJuOnA9ou6J4Fh/gqAui
RCcqv81hl+Uv8BmO5Sikmy+91qx+SvwPm2X9gbkXQKyg5MhWjTqn4SpqG4ywULlc7NSgNspjxZTq
3f6Ns9BEoYrP6egiWEQz4hFfJuCv9TiHtqSz8LKi/EMk7/DGA1kKQP4cfDtZD9kVr1QwivQVYaMg
00koz3ZTAyKqPy1PFKbT1Vm7moy3DF+3utkMie0H/5oFh4FHWmgDeDiL84tuumN7+0IjW59TWcf9
Sd7oRGd86xNzLYVfBhwovXrwqgn8+NVdqZvab8gQHZbwS1eMzmO/k7uwrz6eSnJrJQGg3ijVW741
WMa6Q225h1+Wu5eleOLnf+z3+bd5tgL/Gl4e7o/2bAVJCYlpRPWyy+jVXfIXhFLUNSVJu/RIN2TT
8cytqwT3oW0Vkg6ym2ABZOI8uj5cMZWdVv/sQ2EodYWRThFwPUE6EPp+wFQzy2Uf1ovMXDLXp+oR
V0/O+pqyP2e0gI9DV6r/PiBAdjr6X17Po0O3xejZYnDLYp1DQ2XdZteTuXuOK/20bOPlRBXvcm1V
Hqci+6EKRbHcCNFDUP5TI9nMtv1HTMrfSqxXSURtusOCxe/UF9/k1zFFnjmMjTDn4Yhqbfw+bzXw
FNe3ZPu/Uutxz1qhbNqhGmPh8t1y17cyQ6udM4Qhuz9mRUCVTzEWNbjCjOHnMxkqAnipwiozA2Xd
XCShX8fFQnCPO+DLxq3EqdPiumVhPdmzekYSk+es8TNIFoqn1CNfyk9tkUOyOH4T/kcE9a962Fsz
dht39NWVhWwWbljK/ZbNL7Ah02OA7GtXLlUB4QK7z0QOB8jSHZkFC5LT8KGbeL6zS/trG414VpL5
6mPYFh9VelSfOtQLDiNGbalS4fYENNAzkvyFhttPNdyDe7enCkXUR6gq71JyciV1gKDc7vS8roac
JK34Ob4QXnibWBHrXcyQpc4mo3dVJ8Co+xnI+CAUDXIPld5tnigupwp2geoLUufYz5tvM0DlKimM
EWUDeMbhVJzebJGcFV4AwEaQyCBonldLvc9QJog8WRIq6T2iwSsOaoyOSA7BJ+TGqyUno0/a4Ik8
YKc99uVW31tfJFrUmrYnBR/qbff8qsqsIWn56YEGTl51HZr1oG0y/q8hKvZ6TAV3C6kC2sqGHSu3
784sCGp0du++rCC/AYcofWqpZavxBv1mTS2fFiAZJIDQKRU8cEBp8oj7fOuLmTfG1LI5BMrLO0nA
Pb7oL1R6J7fA5BW7xG+/Vo3QUYkzWsuDE10zxfFMidfBV/19eTYD7PCyi3pIPX9L7EI8BoUB6Pxg
jafpeu49w7FWVkwAK7m7X05Zn36bWYXcFt0Lind32SS/W5IGfidKKLuJyNj/hurMi/z+DmWVcovB
myOlouhN3aGx9HG7mh6gX0AjzNvwuRrF/ne/pf/D6L/UNLaFxLL/rhBxgJnSKAdKlAVxCCMM36Co
q9rLX/lkPtXpSnQfdJ0NJJPBEOU/lkvsMKkZUZppRA4eBvYVJkCqVL6tOKkU3f/I/YPJtonBhGQf
0nH2WPOBFF4QHMfnguDA5MHsCWqMbqJqd5XBvyMlmVY3UyQGNd9kLnAC7I8HZLWS6zaGBUzdQUiM
5a5LrOtNkt4ayNazjeRHhnvzsBzJspWnWQsqL3R9q+pU5FQfttWRwzuVdjthWCT4YrltQWUlCdeR
IwzTOBJpGGOkeBKQFARxELTiOd8HE2Vc0WkR4WboRZYH6dOgOWA/C9pD64lEB4h88lxHHDKQ3fD+
o69stvVej66kfq5kY4nRf+O+VfPKc4YLVdGh63QIc8fIvwWY2/gGU2nnexTqmAHNWpka7tIATrpS
kVtKJqXoWseLOayQGG7cSAqscln51BTiClDH8ZS+ar1p7QtYmpi88UqpZ2GVRk99sBEG0P+9r45M
/5qEF1KLL0s1LKt/UCKqfKcUNm1rPH9iZ77TLotsKyoZ1MKXGjG/sB2oGIoY9W3rqZFrO6gb9cvS
UR1jHFsBTZMlS8txIYW30BGBDDw7XH34kVj2nIGRQ9N+i24RkHAYCTkK+ciSSXFjg6aQ2hiVGsfO
W7bkjysOrqjiHeJeNwAeYtJtYKLMtSjTi4KUKtmXYKP5TDEdTYMrPCHCRkupi/e02wKUvUHsduhD
jHC+Z6kmS6TfzDeE6dfCFXnW+By5S63g4l40EJ+BxnF3c9Ll5NL7yZ+Re8ICbw/8jpaUQlWlwXfN
XKnHnPFYmrF9XmB8N1dytfjJWi+yG9Dq+W/rHz7K/ZAXLjM0uuSu/wPfccDG10QMjX9aVmxDJM9A
qyehwrHMOCyFIrDFa+yXyeFIKhCNGHDVGoVHXqcFZ8IQANkBkqGDNBCT7qjQKLvMmVpzatv4BE3g
Ho5l+sbwD+P+3Cq+kt1qg0VtBK+0SLVRfqRB5ORCof/seS+4PsurO1wqE6N/gDV4INTz18O5E+yv
/xe+lj0yNFhEYbycnp3ztizh2OPQxuatY6ulm6Z2Y59l8+co6BG94YqcW5EfMn5VXem1MzBNoCDE
a8zlhn1xcYIuCvTVQMx+hFFtcHzuDtbgpuqzxWuoF7SLWIvHrdTre0IOWM3r87lniZEtODJ+jx0q
j69QNB8P2n7kxhBijqMgc8ulL7WsWuRrNJ3DlM2f3azP0uGh5CJsQQSYcGBdJLnxskNiIw623ynp
xLMecJEZXr5LYWGc+lc44XA2oRz17l1a/9sOJLFT1kwPzafFw7TuGrv5KW1VGWDT5J+AgOqUDS7n
IXj56CUEDOR4fXuYX0lC7XAqZI8XvRHYmx/fZ+3/DXxCtEnARvUYH2OduyyXh+UCNQdOMKDsZp9P
5dveseizkYIcOTjD7juYIIGFMns6ehDwcaG8cUQGSIT64WRC3Me5DmKsYRsuk7/2BrtwNxlz+QsX
md6ePuAKIz2IsDoSBsTSNbinsCSL2dy2Pi0U5JUlChkRB5u2E2pWRHS7g6OvhLhptNuQPr0CRjwE
OgrhMVdIT7p9Sb6mT90jo03r6S3Y8dvZuVTzRsNgjDYG7xqJk9dFaen6AuETUeKm5qgKv6A8h34/
qQTHLkBCp+66EkdanLe3LYNiRildCeuNxf7mDE8ey85gT54hgjTWi4L1b7z5gxMAWRx1jOw6wId+
34gLNmAI5Tw/2jybH/4828ROzuzdEm3e8y95c4kgSPUqy50/pzpnNss5Nu6+YpAnjRtiCeU3lX1U
q0uuYkIb5D840+XilamCUuvKlaFQUHk0VrIUgzGzUc6cNsXMujDmwsQog6gZ1zrty8dXTMf+rVuj
aNKTj5eHKXs7VoESCXM+KoZpRU6UkJx//oQpC7ziJCGMGG7jmnzEx39uOyHJJoLcqSu1dCcKJLX2
PFdIrJgLUWyU/Qc6v1gV8WQ9EjBl1xK0pKkOI/l41Os8+mp+E9HhvftwvskAP83H6NfvK6FwY6xq
A6Sm6Yf1ygZNJqxOmvW8+IkVBbWwLsG2q8/N+ky1HSG1H4v3PEuWngIL56IiuM5oZdtdPEEOkcts
tHr76cz2fzRJHHhJkkRyjjhSqkl8tES1G9+zNsR+ec8OseL6LiWFH3E0lxSnjwNgsuKk2fz8qVDC
INJ6R3zL7Ny3oTaAGz8D85Vhs1Fx3hje3GWDpWGkplsdpVdM38XJH4MoobdXfRnUWgp2J7CVHa4U
p1r3LowZbTW7AUe9CmFcI1/pqbCa0EA1B4ED+Pr9hqCNZ9AuLsQ/hkxbjlXQwYITo0c79Bp8R+0D
ShgeY39cJeXmzerpz88Que3LBvaaz+SH8NXGFfDlz2fvMAd4aF7Se6va+AB97BdpNm6rxNj4WlBj
QIngF8v+aQCuYiamuEBBiPlyH7+lw7/ElhMgaAU//44Nz3ZczCteLJA8nnlovNwVdNaRZUXgyKMj
3vIfduR7FnILDhODg6vJ6fMrIenDsRvpuMPT+VagvxMf1s8S95moDFUPfq7xC8oAv3wg+XvD0Ygj
z9jDa1yDfqj9KgbXGowAgpXCzoBGZ70s3sDBsRG8FmheGvFfNIFAV+/cl9rXRIQmWQLPmWw9Iw4g
BriOYpvHySIDqcv4sGaam2kdliqUM3InEaI4UzXO1yB+Mp+6MIhDZjmh7u3Kf4DWiFPqyPKPGDAc
p2lQWWWRY7iXcPe6V2f2RpUP+4T2qWH+IiA7G3Y4/+YMuR2lBeKJuKKTBEA+NrC8FsEjbyrmCh+l
ajvsagavxdSqlocfvSxr1k3D84vRcuFFs68JY9wZpYolbaSUsv3GWM+82Pygfp18IV5Xv8lUSBlx
m9M7X2wvHPE3su7v4cL3gd+fTNEes/3PbKdOU8O3dZJk7wmv4xA4CGRgxh8Exm4SQEJ2Ix2oeHlf
SY/rizzT4CT19UzCkLJ0tXAjhn+bPCVzMSEfeupTnsWIQ9Gqnx9ps1z5iqy9ubliC3whqk8TmXb7
2ii9YZ3M/WvgmdxLva+GeR+NWn6FZ94QMcnAmOU8zsgkUdB0+2qWiZe4Jkv3Dol/fEGO0t1UKEHs
pK+8VhlJo2Zdgo2Vr15vszc0zUqzmZXlK5+/leGkWOrbVeYRaMghvx6Df6NHDADcm6rFfPBixiyC
KZIz6plzdLp0/tiqRtDW4TMQB8Zymsv36yRBf/xdy5CFDqMAP8tn1c+VYKsOd6L9nFRI3DisX2H8
BXxBsy6EOeCdlY3DS/6yA/0Evtr7Jsw68vX64Cnt+YJtAxS+Pv3fpCEch6fBfjKrWgtnlvYl3vCu
2JHkm5L0AJRo+mGj2zd5QMRwaxy6LD/u25hL0jKJ7LpOmmVUjwaxi3k2x1r+/JwqWJ5AT28GDZr9
0c0mAhHQhc/hxBI5xIgVvf16wzpXMmKIx+ssBVPJp9tu1NOOh1ysTMdrIkvzOSZn53AzFqK4McYC
XMqK4hwP8x7lBg+Op5WVjCZZ4dSt9cJ0vOQv6RyCiUQirRv4esB9NEoB9GNV5F5EnkY0FRBmzCal
fdD2LxIRAGcYSMAnJwgMTBFJeote/5/PwcllfDEOCq6fA+vQ70CWYZK3ZbPD/R1/70nke+70fU1O
H8lQ2+BuDudEG24YlvEXtVmfPNZsFKhhXhvzXlHJ/xmIBdbhyrPUqy7uWA8v+blnePyZQNYoqjKr
+oe5P522VPC8jqYI9HZZHaHJc7BpgsZ4SnY9nOMHzZeJAK+nRsELVy63ttl9wLbQG39ToXRtWROK
RYIXccsPv+d4mRj+M5T7hEcvuRCpehJkagKYsljWycbIAC8fRKnXHELkjIAmj4tTgpOBqE/ro+k5
xL+lkxaLnXuuGD6u0dwFC34l9jJyow8JJ3XheHIx2tnizEOe7ltnPxeQUKYH69J6ghrnH+1r3twh
Aca3zRVzyYxlBgDqJxwCMvYkzIgTZ36WNh6BLeq9xGeNv598sHOKxM0+epYzHcocQCzXrAs8T/XA
YUqHPrX6UvdeeCiEhkbmAQExY5OcsPX9F70AmxHPctgupu8BfHKj36LVEyWhS55ZtZSQiIw3adb9
7t9by/C4uaJsoTzDwLDBKAXVyEFf49T4ShWYDHlc8WL5WLe2DhFT0ePpg/BSlL6zDYSSCegVL2Bm
7fGDH2MEbOC1xaJRKKHzcNPFHH2lltFd5EEeOqVWf9bw4K6ANLFlO//zMOYl65FG2q6NAu3Mk7x9
hUp9Xn+XMpE0GFq76S8ZnBu4fyAHa7FDErToQdj3fBL/gja7VpgvQqvaZEI+rtpzTL04+gXZ4C4a
2rkroAcZw116L3AAT/6dqsd4GGy6aaqtPaRxj9cB4uGwynYSm64e6u9Efj0hrSf4Viy+lbYBi0pl
Y3Dq2GS8Ydq1uJOHt/nbNIcHEvt/UxOWpCQ3gL4Simhr+CNh/ye00kyZievRFLTekDYlIngYx/hE
frXtX4x2Ym84cEo4x510Qi7mM0vRGmrMoj12ujsRvQ+BLw7dVNWmvok4R4BUz+q2iY9r1bMKLd5w
v2fq19gs6I2TVoUrJEMtr01fBkEfmh2FULvbv5KR3ojBx4PPTscZKmU7rU0fUbr5EZ1bssMThN2y
qJAIh9QmCabZL4cMYhU+0voJvaPQqATbpIhmA9NE7v2QQevqiNqKcF834qk+D+RKjEkBmt+e2geq
kXZ6QPscKqdxzHHECsLHbNWcYcWpN/sb8nJj36zqEO8UJQsk4EpcFAqA40BaDnnFcmAYygz1NFnr
+1O93DDSq/QNoCV9i7Mi8YZFRG0MWWDaK1DsqiXqBY5fI53OKDXjo+S2fIDsYyp5MrAkTj8CQIb3
B/guF0Uxo5c/UMN6Wd+m7LUREvoXZIheC8X/K/NpEzBRZac+hCggzmfFd2RFLW40JmROdNJK5a/h
F1bQnxOa5/+x98FCIevXUTzHMwlDHd/AExU+8+FQNW8NlVXy+WeHzAK46hA4Ccdcnut+s0E5VVsd
tTk419cDQeVq+Th0cLC2sdW/+DA/7V7W8Di4m18Y5DO0P4U4yPpqYMlNHYZW+wwXVL5tjZoJBp5c
3AgHFX00hcofLvqVBcBRFeKPrw2rGt4PLCNQTQZ1Fi+Mv3De5UjZjA4Sj93NPhko1X4pzWARHfaX
1rzLqPDWwy9V5fGM6/OIw0Hu3+ao6R2y92beKSnlAw1giAkrvRFMjjY/OJbaNgqgliGOhsLIA4GZ
TU1ly1XQaVY0xQLgsU7YnHW+hGTgshCQTSsJeqCLef4cu5GUzax4D0Ace2Zt46qHC3o6wGpASZ8A
3RPF1JKALrGUVmtLXglo1GK+OVYIaJnwyqq1Zu7pgpjjsmSMjIMi8Ka56M+NO1UUH6OGH0N04SMe
DVhLyJfGVk5w3tL+5jwJRSA0zMz802ULtCJIC3O0cl7ehxpnUD9ahySFKLrrr6vO4T5aBKlgDAJo
QSRequ253est3caJ9tvMRGl8lykWsmE+qi5TmvRtEO4GoeSKgOgQa8M/VmDBNSlGGafkyND/OlPM
v1fhCj8j5CtRhJ3E9++/yp66JRFYeTfSZsjMzpa4iRJU5OjUaC0OXBDktsyBgJjOcQVDoGILPZ1y
UkHBBY/aHcNvSX1HRiGCu62oRV1WmMx4uygpX/Es9aNIjR7BDK6YbXg0nLoUSh7SdM5ogZ1rqzG7
O9QWGwKpeId5+02ZAJIq7DaYunn6EDWGrcGBfymOJYjaCMVYu79MIsOGZ5qCax7+vL7ydt29gyOM
bYLn2otGWHuzREn4Y5GOfoCPJSBn0ba99OXhvHvap/M1ERvsE5pyOqpAbfd5NMta2qoN1OFboic8
hsoo6scVWjgYP3AUEeO7HulM3ipV6dFc703Q+aQkj7rlKNkZ7jUYzsBvuxvw3X0IZfTCDj772S14
enPKO0wQENS9rj0DDHtf0cZ7yilWyh+m7JcuxhjWPFOOBn6N4I3RVRJu2YvsM3qBZ5vGwizKwaEM
cRNYSswmm3gQlu9FQIeI+v16rurGxxEo8/qsuB9eE2cL3nLSjcsZXsdrv2wUgbSm0neVBEY86iCW
zcTrlVGqJ6dmu0s5sAv+OCn8cAYY8L0x8gusV/UoMK3pir74cy6hUNVbWAL//nbvQbfupQQkDbPN
6UAtBpkQQiMxyMZeXmBugml6liqNaEGb4CyhY2HxPAAh3NTV31U97UfJIDtF/AHYOirK91YU/Kqt
+8lzlaqBlDF4c6ongfLfJmMk2ghlfEmTdiSGvMbkRMRildaI5PkTVYH+Lfvp/Ip5Yu21z9CFo8eV
KdyDp1y5jMe0vWsgiRU5ZPMc2nH22m2AIABnwi997U2bwWZPFdVzPyQg/Xy+1bNpGbHBihxXTqL0
r0dPQZAmyaPOt5l1ZPQITQW7NcPnAGZuNpn0FoYYWuiRZnp9OCVNbuUdIp9P64aG7lFgE+xt8HqD
inqOEmHoeyzBcW3wctoW68amdKDYy8jPkxBshS0xRyIyHdW0z1MInYVSVW0adIM+13om34xZr5yX
S5PHg++NmiXwDGODnDbB74U2o943umE8zCsp2ijNQWo37/mAGVaDWoQs7QuVZc2NU0cQxdVJ2bKB
AQqEHy6Iej81nz6bDFSQrMzC3OFfH5d13Krvw25oyUCu9rlfSC8eGbT6mm2nQ3oinH3NbklOALL0
cqQQ9sKBfGKt1hINQT1JEMYqv5On1/PlBn7sMKtZL4/3fKEy52YT5EiHu53yBQzfBbY6ZVvRPqAG
+0h5KDJTpTdAL5s7pNoodw55qKrbJ8geN2afctSXnNYokTH0ox+/GvNtPmx3reuy9ovd4xBvTdeZ
gVLM/U47k+vopJH2bP4lqPNFB3glR9ZSXrp3cHsBpmOcZrhiICqYG9jPbFS4cvTgEg/x+HOgnioC
Zx2T8q4BsnwlE7jM8Nl1sd4Ge5IgtiDxuZmlgfGuJ6C/m/JP1Ju0A8NeqSpbJh/JWyJZcOSbLtMg
TiOBmW9V7HXSg0oeDHvbLi0R73t7ezp16sJAw4smw7k59oW9gTSLA9kxERZux7OmF3VGeWZPVmVt
BbkYZOz3v99v71gFmfjOHYEvFN/D/Ek/jq0CIBRS8wafIw9c4kkQ5NHSs6LvYhCDia9Y3j6Ux75B
9pB8BvAmxtexAg2xEwPKTvXXoCG6MQkE7iHEJxqbqkclOaxkzsmkDA5Bay0Jdhw4bDatcXC4phDe
NVmCVeG9IsIJxUuZDn4BVSnKUZpHPPAb4tOzxj/9rHoIjJe8jTQNXTUrpaj4f/faSI5SUG8ig4e4
LVN4hbpAmSCkY4kEYOWfVduJJ8el+BKoclVM3GA0MF9sub0WCxVI5WQLHwKdbtHMpkere+Dcc9Py
qz/zvPFGqdYk3OsxdBk+5xjSQhx6OTLWDZtmay+5T/c5N6OTPm5dSEaykFEvuy2Ft2OaByE4qQm1
4QmcNIz/i+lwxvK5MdDnpkn/8+dd+1RL7aPtZlI78FlL6ZWwv073bKNJPbYvqKxmHuXZzkHSuZyp
0q+yUsackrRP3CMQv7B+7t6r3gsXZcGDyqnSyyJ7CdzuYoavokTWiNJjjGzFfM86Ue02jERhvN/7
3r1QJ0Xz/tlzxYCcmecq8Q8LWK8wRRp9tfFWB0RuoPaXNkhGmgA/Z8cHolUDKXLav9OFrp8Z57Y+
ZOx5UqcjJXk/zBobt8VbrLwyO4PA70rQNKe8yde52rIgaWMfOLxBgWLCG500IoWE19igk587gp5Q
UjPgDwt16IpjCU+bVaomvdCvxaecQkSOT2L5nGb2zWkGJPqMCH8h31S3Y3s34gTOSM4HLQg3xomu
vQJXcCdJstqaMTR7eaZ88nNIhXf1Sblps24cRfQGKyV9z03KomG8/kY274xau86tOWFqQOBEZfbS
hTpEtXvGgQ2gdqnq+nTSjsH4rjn5M2UnAP2lKqwl+YTOIUNiSZzw8NdLeIpOOamrqmvRtgG78Oag
7KhqOJpvbBRhubvRH+KMj9t7vcMKKCzb0NIShWr5xwtfEhOpJx8iA7LiJy57xMdnIv/WzG8wrkxy
ZYHKtUtFEJvYVV0FTgJMja3qRMvYZ8mhhgrcGNliqEzgyEJLMPm+KByMiWHyPqXjwQvfQNIsm4af
PfxSl96wjwqsSrCTjXQFMkg+tqu14iMw7AR7XvQvJv5KS21oZskeTT5EVE3ORw4xH64KrbNhnF7+
m4VBN6lKj+uUTx6kWFjNNeiYzk0dFVvpaGfKgBmDJH0EnzrzW2foIdroFYIWh/wHW9aY+IijoP3Q
cCvw88a/26UNm2Lfd5/4qbxsCTQjqOJpOMxvSirzfkwXz8xL0jITUmB+r2CZB14rMYARf2Zr3EwC
NUwmMyLtX4l7ZWpAUWaiv6S7IAd9JTOej/siWr/8qdSE0COKBg8mSK/qHnJ5+QP4vDt2N3J5Irrc
nMRslpoAGwmwtpVRSxGutdkx5BznxQMvMDK1IlYl+faXKsVANfgR73cOOcPObswPHEFhBz0OzvoC
VoCB7eeKrsU0dsM9cK1fQeeIkGbeygrQ2Ozg9dTFSnxKgjUEcbYQA6v9+YLwNSuXnQFaKrajxG95
Css7W62sfEFp9qG8gKrS2QMWcI9+DcQHZetsChv5Jf7sO17TdFVubRQe78oj7M6Vs2B9+v89XtAL
Kfvuzs59g50YWNvjy4pvNKlND/PiIyAp5t7OhWgbTBenLVhw2/+bWp2PlRCu6C/C9ww0dmQaaz7T
qrR0kVRWGDzyulzEfvo5yjvMfq3gEw8BiWRc7A11zo9oZVnlJJ08oSmwzrocBD8iig+4/7GGiuNN
yVawu83MvXw89Cbk3VPOzdwIIx87RyUES7xrRDuX3aLutkNmq0h2CcLpxU4B3DMwUCQauoq1uyfk
kVc2sLr3NHV2a5T66QF5sWp5lxv6k5SHbiEuTB3KglqGHKcEp57Mriu8AfEGQWLaQ4+HHIktiZEy
TgSPQZFp2j//zhnrKQEWWvV2/q1ef9j7tcLdEhKpWIq/XOfO3ohqqL4ctlRCWTvd1yPNsD4c+Xya
uwJcBrPbwsjrBKhcZKI7SNn0zJ2Bo+pGFJHFnCeEYkD6G1KaWVZqzRstfy4A2aFfl/FlXO/07lFv
XdTb6Fy5cPuPgYj2bbZ3FZ4v1L0o0fplXQ0yycP8LldRihYfV+FMZep7tKHt1Lxw9Kp+UQDdP0oW
O2+MQszGah13XJtovTh62/yjklWE1S/UKP2auRyMeIFWd+mjovff+pH4MXXwas9/TAFZMyB3mjnq
aBaGlEwcR1zakWdcbWLd7aLuppI15zfsOKS+8KZTVrDckdDK+wL7Eqvd8dzLE3UiZbgPHcezcWU+
hhuuBfSIQtFNSCl30gt8PHzC2Zh7gI69cxMOjZR2foRjlcc1cQp/GyIc3TTCWp0so+eEElV4C7UB
yrwttCIsqwrfv+Yqj7vXw8ae0NrNowWyH9HOtbeCVSIxErgzZ4JPvZAufqZJv/GnyTW5XvEbh59Z
71XK/ECT00+hqehi5MNGguIAPs+hkS32l52V2KFqY5IaB2VcdJ0I2iVdSbC94u1BofLSTlyRZ0zK
wSPErq6mOAPlv5vRGR+vZs5OI6rYaDgMPRi1YkfyJ/QOxUQXxO7QUyMyvqBMUTgFc3ud9OgLHgys
TQJ+bYlPSgG12qVeTLlF8a4XY+T2Uuj2yYkqxhhIW0d/7UCljyvsaQ4E+rfj+n/5qT9pL9uUa9Q3
fNc8nwzqXDxfezBrJ175ufkEkgE8PFzK5PpieiwgxxRRZlhnP26xt34HN39lJRgz0twJcirdGVCv
lHBS6dhbPhT9p/xoGxyOsEHhEYSPT7Bj8Q534BFAzj+xNQCYNRqUmRyGQt6PAwHw6+dWHMujyVGd
/SEXeqd02JnmzYSgpB/RUiK7cwrL1RjBY/IQr5JfZXxRT82xqGO9Mk8rSqLahxYrQjkiszgYgr8o
gzQPH/yMJkGcKb4bpj+NsZCYYVbUAYMvdgzwrCzf2vBuiqxFlExWVL0KcGfrGiKt6+OujuzegmtT
qtZFa2BU0YVvPS23fpusaFLTHuyh7p2UCjI9upss1WBAXzeIf6bNoMUb4aGUKGzX52V9/zESnD/7
J9uRP+VyAeNwC3cir1Y8F5Wtn00+gMHzWMO5aZI3wKEVaBuKvd4Q73ysFcvLWQPKxpW5AMiKX/4o
0Ugravlsbwzw/8d42096FJqFwCSP72qhld7GA66F4jpYdFUAPlQ0JFo6OAB5XG5BVmVnObebojcq
b4EYCPz/DqgveM5mUGEY6DyBBum3CJtmL5AHlD6GUJirVDhTv/T5Mtyv4Op3MZbYUr4K77uc3G2a
DRew6c0tg6b+g5LcT2LTCszWWlLjqTKbncsvRCe93WPvqocHCUJBNTDw9Pf9IFNAWEFoGumxqGyb
8HzN9ULq5CWwVOtS+Nq+0JhH2PEf/DET9uERlIBTDozBmjGpTaPcYwWoGz41hFJ+67RjeVtscXMy
f5vImrBVXDqD73bSVfv2GvqBADPj1OtSjdJQk/sZfpqdNCLHZ1zAb00PsGa/VX9rlHrGkNBXPmMl
8IgDQpsLRmQWvXboOTuOTHeqFwZbdETZnyd/IHDsXXh9FrT4fnppt2P5xjyFw2IIZUSKMri+6occ
fy6kL2mn9wCl8hOwi8j53GtDVG6zY3JGLCpnHh9dSypbQEDAG6BxsFL6fUT0o4E8n708azuMH43H
0wpbxtF6jbwXtWiy/efRE8EN2kuM8SqxxNKpRhamQlP4iyUglaUy+dRQzBceJEqs6RhQZ7nlUMBF
7XiOXcf4JF9Ky9mp4cEb4m5Dp3mTduy/6A1EHq2L83XwIbecFDf4vG/G57n/gJw/Q+qBTyGkyd+d
9DU1iKE9z0X9q2Yiu8KdIRi8g/xlnO6zGVCz57PslK6uEi1hJgSqSo7ba7if8iu2b9PVB9r17Rh0
mEXvAg06S8tqkzsw2IMOLl7q2lhvxQi7XygxkyGZ5IbQggS6dpi8dJtaR6Z7SN+8vCBAxF4axNrj
m66yXnCMjYWjvX3Vx5jO7aUOnAfAd9VcZjYfuJxNFb7J4YOL4JVZ96n5s65N5ke3BZfJIYBbG/P7
xUi2hVEyKu6qjmI+gEPurA6syXUFRSrefy7wsVSyQtKMQ760goFikrrDCB0m4vHLFti8vni+s0AU
jpor62qoie16Oit4j1uadzJT0598I68vjvtEpBsj3HNW9ZQX7D7+WDhqiE0R1DGgDD5rniatjn33
dmZ3qHEYmr68ldCe/rEqPBgZfogC28WrvwNj53ncaPRpjxbwjZ4JiFpByeT9xVcmx0Y+BIMSzHuS
aBLY5CeUZSLcgnLA3ARv4usvgkmmV+lBLr2DCjo1zOWwU1+OMYbOmhS4w/3+24L17TJp6y1Ndkwe
QLwaUNMIiN/cwUY1gwHjYmHkoJS1IZDewxQiRlmfj0b74y9FbWmNeDR591RtFeo7bAd94wTACwSt
fzcQ/xWEfHujkkA/nXrosIOd/vkGe+EyoQ0W0EzxpPGpT685qN5j4IlUGgcE7W0Cst7c0aQJnRtV
JlGVOjxGoWyX4q6wlQMZ30G8to05VUzZaJRSOIpFIffSD5R4IsVdTUD6wignkhrAmCbk86kF9e3f
k+aBGncOeFhLro/e63U4MhnXO2w2mOWzbDZc3PA9TtLHZUF2XZufkLoZ4Zd7G5jo4VpwZrtouSHJ
+RTx3fGmXJGjEx4DmJrBQ1UmS5XK2AWBffBMjgabY0ZA4mes4js9VuYm5U3D/j1XzrUIrkYwGIay
B4yPX94MSTqy+uVkzEPugvQuTvj41jCpfjlNv5valFIGAOdDoS3pl4s5hPTdNsit+l+712w6Eixd
Z523icdpUedSBMXQkaoWSdX0oha08qVK8y9mFFzDSaIzl+97Xv3n6BbPse9Kb265uKQ5L+Jr3j0P
vpm8g/qLIJFri2sCy+jOhndYw11EZNQirPuK85CtgaSJDdxCHDXfVW8w5+YG1GhN0YE0/obFuHPL
yV3IBGRzRhofhdHMVJdiTAUqULO6SCVD9SQOsZ3cq3W4JsHNUoh60SbUPXzePxoe+qS1XThSL64V
ebTXXxYVTKvzD4VmjutSd17qqKBvUOw4PqF0af/qiNi7EYmYfuFHHP2PFkQeJoHr0xuisftPWBN1
s4/0beN34lw68nOB90nbPtGkkfImI1BaSsyA2dnde3aaXsHJKBc6uEMGbHRfTQIrnkBuyECrqWg+
pG3IBEffC+QsZa7RlF8MeVhmLAWWfVHSKk3pgJrWLiIRerlj3HdtgUPqs2CT1KpIVeEDAZv9GOfv
IS8zZy5gDp0qL/3d4m8IGQm9zSIy4XR6ih2BN8N+v3m6yXHMqJPuo8neEjbNw9RLIJl78BZAtiaP
P70Tr9Q0jOvuLa0xtnSL552ncVWeEGkEiheKAj/xu9mBqn6KYwyNeVJ9pmsdrv82TFwSsxOrybH8
i7J/+A4syTQ2NsTpj23U7ohZOsFQoJvgRoVlznQwA4w3m6p8BIvOfbDc5QevmkmvJez7uJ2HYvX2
PrvzBoIOLAeNZMe01dDtT6naebK5QBIAC6Qp+iwWfrYVyjagZ1jl9pAxN99J29YwqcbTnXg5yV8T
tacpVXyugFB8/5PP5Fv/2j0rD6sT59HdkW/0yyPR2AD0oRHlY2H65gteWG4mX1SHTQjV1/f5NQ1T
XN0W5A8L3O6l576Mj95jY9DOjAGchhrQEwSydqEuuhk+TIy5RXZngsXdcDxYTodS1thq6qkwtcL1
OKDUHzX+ZDQam47oVlL1ZBPCyOujNWJP6s5EqBwG4wDoLC7Ncr890KxkP+2tCtSvIQKGr6sl93Yu
0kZSHmvbJxHBHDuE79Zw1dbExeNltqJADz5EiypNmvoQd6Bj4iIm9h/8dvf40ZxNqqHGx4rFOW1M
I9xUXBNWb/jv+Y0nZSQr3pCPw+3XvHvgt+TNmlbMHvZTlceuIFC/notU+Rxvblg21zLoSt1KlGdI
TcYTh4Qa2y/Oz0VqSHRzOpH9wuLIkEZsUHeG/XHi8cZWMo8VSRx1wHyoktV3ODUe9ve7xEmOb3Pf
ZSnl5DsEJXuptfVUO8Hd518Qx98vmkk9QFlekKZvA4lSJk4J8BW9QVTTwlKOQW0ggo+43spinmv7
bC7QRe0xMLxELNOY7/0ULjVn28zJzbPCrSkdOsY1OkwJZcSDpGWDMzwuVzRW0Owj/VQYVDYeWgve
ZkLKZjEu5zs9Qzkv4XAWhWwV9mItRQRujQ2gmQ032aED1FPUAdoO9+EW7TqajDzmJHA1khOx5mN/
7EaeorVIykpWZGC8PRT9NT5+Wc2En5XA0eTxfqJY6cRrukk3gHEvHQ8zdPipTYiv2kLZ4hB7Fnpw
gvUc0WmR6/FHdH0gMIgD/Zztp+k9UljQcd/vcE8vS1wcGHatw/O9UWIs6JuMH4KOJFXC3LsJ8+/x
8nQpL0ZLXlWEIqklwacNuBYr5nMRL7RXVpVW4eYznG556oj/UqxEPIQ2BtrVQbfpkBdNqwBapIz3
Gk7xlXFu2z3V8kCGlafplRnCmjKiKufAOyaxrDbcx/wdUGVaaF2FBJpDuvr2BtG5GUtWNieiGtE7
/qmEeoxWekEdc0gM3wB68z0dYXvppM+RgHj1WcfKyO8pCctjLUFdgP5KEq7KORDO5teFqR10lSDo
Fs75RUbu+gBw2ywem9iWFM/LTQnUsaub5uIayLgbO9XBT4IepZgB+i92kHD2fmfxlxcELaGEFvhr
ED5kecGTHGSnTghlMVodCwG82GHjp1ECrtR/GZztaKIcDSA//vfiBQJr/0l5YhPjkeQJDPw8vk/M
DWQIssr9mrqdMV4L7M39DXR6eME8U88FYACpe/SPsXweyTwPMy5fS7OeVYNC3CVR5ywmUAEymWl2
3YehovoNoWY0CqpYZW9wTPOT+OEaS/FHF0DeydwPYOR7tE/s35rDRiXPLFPEyjOQhMBsUBrsnned
EhmH2P6l8nrbqswXgTUDirMCmSrBH7VUFRrd3qByOZMMbr8Rz0dZFkgrCz1DGTOMY+gET7fq1fLu
qPMFxKA1Hcz8LMLbvOsUHztJmFGCmzrkk4n1Svn8XbN/ShoiD6Z5HXJtge3odw3zRYz4tCNDUybD
tQZY0PVTYy092F0PulQxn7QlScGinTsvlsPDKlLR91IHXoqwLyxavIOsGXzx1u95G8flRzjROnGn
i/09aY7W3mkCDJxi2NF6AvYIBTdlYIcz9RU95wy6pZl7Hw5rMk07bWzxDpueRensxVFhgmtvZKI2
VzZ61tNwIaLl14WOogTDwTI2eeMMKlveeUB+k+Rywajj5wOBC5KSR4C60hWf2K566PGb9xVkzQRS
5D8CiAj4xHyxyhFAfLygyPZxrNR6w6FSFS6Xseswa61NgOJx2Id0hyii3HaNem/rGbPJ/fgEvCmk
PmCSimzsDhyt1ZM706oyWpfD9ru24ViUSvkI4Xsy4f+PwLDU7fQDvdUFIRFAyfXUh7nAEyk4bRtW
Cou/LAOqkR4F3dAruTGNcjasjjM8lXuprZ5iyb0NehLaJGWUR9QXQoSzTQDYk4ayT7EGGZHgC/oH
v2wQ7uiBSdR3JAHzhg0Zz07ErBXNb4UTdISFitdBMqMgR3sOh+WHiq3ILgqXwNdYwkeG27+sf4CO
oRiEmxjo9BJDzbb6/DPBo7dSS4AVlNc3loa8byqeC2mgtsptZ6M1Hpwh5bd6gFQny595RkdACmSs
Nkyaf6f7jUrzU2Kv/ebkLTRHbUs2TEJX7kBMl77SlVxRqACcVD/0OC1i+oHzrUjX0RiK+IA/+5aO
lzEWxMiFbpPiHH9RwQWFfkfvjFzJRh470pmZe54bihy7Fpa0PPv1xOM/ytLgMEdWcQYv83eIKlMj
lyOL+Vv1aBA1DFIzc0LH7fz+D4eHL1rm/rAmgBbwSCUEH0rFr6Wm2OZKqKGJ5JIeiOQldAP5n15N
g1c1ALtdL/4MGo3iNxO5+8QGaaWoiQet0rLEJzy8INF6WE0MpZZ24pZySI3FtBojyJxHMkdXEfPw
2qQatR/xIT/DTiiYfqn6J5dctaJ3DyR4eLZKymCQEQUfRMYk3dHhdr5WxkaFvh4IweiLLqaDWhwd
0YbGUDLeNJd6/SIMGuJ0sNKTLco9vidmPJ7AD/eWuuQVNvZssMKhJAv3bt/hV+SU3HPMoVxZS89S
WlRJEtKAH781RS7NTvwtaMvQZnsEgFhJHkzudPL0R2Eux3TmQNgrE4ACubtAgpf6Vl5PbJoT2tjw
P0yPa1DyPN4cgHux16+P+rYfu324yd3Gf8Pn7E0txR+qZ1jKTtqY307vmhhIOHBCs/dP4mgTT3qX
hXCki0BNxF7gFb11+ZbqSVSz/QTOqYL0KRLWOMmKbcJrhEUaZwOYahqHRf/Hf/lPZYSfQGodDi2p
KoSL0lIG2scqP8GKgOpUzSbHVQR+oKyCSkJiYBcvPjQO2klA7szq+1XdNvJYmvmuT/3dzp9kRFCt
Cdd2YYLKbRIQtopxnp4pRshoV5beLpNg19V0ywecMeCHuTNweex1p553IBqVkf/6K/304MD+pE10
/E4DiOPKLDUSj5PBY3/ZZnawfupvaEbt8OqWH1cTxZAzKxaI6XkMRP2fs9lKKYRhEot6xBQqrXMa
3qZh/GaVf7OVLAGXb2+q8jvhMvRoHBEaoOasAyErWObAee465yIQk2Ue1tCZ4ypJJ3DS76DkqJE7
rEXYxO/KDjfXF6yuY1d/15KkLxaUbW3qQxRtjHNYg7U3mi2N8y6RYj0LJlwZ2M+TePiPIgV4mKse
G6gnsGM/IckWhnKNa588y7MC1/z1hN52d3+eCP+M68Xp0fnPEMJCRlWkCFCbXwZXGhWTEAKSvVcS
saap6hHm1hA7ctU2PWRP2ep4zU4fJQtxceRv8fSWP9Ljyk73jebZeiqBSdgTfEtCEstJQYQupqOQ
yP0/oJtZknMqEy4tNmL8pGZeIRem6phWsO3WfVwIfIytH6/5frRAffr1l7sJS6hszVtbHKOvVCz5
nDysxx9+zgXPpoCsGdcLp/1JM30FDjvjivyz5F3TRFLXfORHexTYQMVNy5upcOwNtGh/bAZZ/Obf
Sjx9jud6LNOdyEKqpEkEgk3jBhCwfyelBbOFtR4vVBJSTp8gJChYOM2/nUAPeN1GAXAAVvfMBoYA
rk+UVySPBoj8R1b5BZ7aNulDuEYEXKKeTx1K+YIdbseqXpB6xkSkQSqW1ZCJTn7GjgXwVHzh5J2x
hL+E49BdQ7z6IuU5H2jS9OCxlY/Q4g3MLif9o5XC+bscZ7Y+/1393uR3q3xbo3k9CdYrHiQGly+J
A/41v02zQ40zBAfwZr8XnG7lMgjJm+mnVIdcAFcHLRp3KatrqZmcJCqSm/NiKkMNWFyEZeVRdi0p
JyuIBC9m/sn5R7EeFTJc8RzgLFzXLERqw/TmcunrNMzrSpuQeFGEZl9dDJ+P9Y5ge0kySzAzUP4D
1UxaVnSxqihICD2z3ns4gmJUNZeIjv56hC5NeyXIlLImS+9EMe8+pX4+aB6i0RoPvv/ymLQNbw33
oUwRAqvhnc0vBoVCdCHzPskCtnmbJ2rEVaa2MEof8Wl/02ZDOtkgVmJRo9D3Ey+Y3ywUbyfIXIwv
N6YpbkiAVRvZyQZlFkZ2TH68AstbHbYyjW0YcORmYDi37bdD7A5MFL5NhdTqAd7mDQmA30gWSWzF
OD1tfq3Xbq/LpbqajurNLYKllQT5UT31VHLHjP1GAslTHH74OP1CYEVy90/yCTf4+A5tryaT9pWI
/NWHKxO0+0zNSRkcP/e/ht7FQAbco5p+PcHXd1k9GevBvmXr+cNyduMJplg3cpZUAM6Q70qGPGKq
J0Yp3SfleyEAY4gLwy+ngKPIux26DJwpquvwlOJ7c9jwPTTIMdoo9rKmqRVSndixF/1zZk88wT7r
dMLmYJUaie6PAhHGutZrDdNOi00W/LNA01n68Ypel6Jem+DgWjxhfkhJ67oxS91+486bdV0ieki1
g5Y8W9Qj/wC4sfGbcwUhIL0XMzu5knPss+QrnZwsdAkcbdva9cf0BurkOQneOmn9BpPRt9nIi11T
cN6cEDDS2UZbfBC5SHly93sVWHtK5bT1Gb4H4kR+o2SAm75/eVOtEDrC7zkKMQ0jXLMy5y5hgh9O
8rni5Azmpe62XNlwi4w9FXl4yv09hwCI5tbKdfl2AlpHx5qrNuX7kQoutQIA+q1Nfw6GkhHAG1rF
Qs0WTLZZvM4MROoVJxzMt2EFTDlyYl2xhTeYwgO8WmUfIYzaaHt87Exi9yzZCCkx6mTeByqZsCZ4
3o4LrfyTgVKTef6fkTHwQ2+XyWUT1h6QgvF52JjrYe/cm5B2fk7KH5K0rikldoFi5SZ2DShjQxoq
GAGTWdzSCUIkEEtmT9o+pLayIYdtSvHnHB1mITsCInf39wC/CM8rML9LRailypZ/t8xeBDEcya9n
KutEKQlJomSHbsyGsC6CxZ+UgBlcBti0RSnN7sGU8D+47o4GNlR0Yg+tJZojDIKR7K6y++ptNoEb
X4FYIOn9sUD/662KhQzWB4yUCueK84pSF6LEV/edy6scNrXezq5EPgrF7G8GsvR293A4SiBp3bTW
EYJBRsfvbMKeW3my2KHIMXl9BVfY7vutWyfyWiOmzJ3c3YHVGJqJseqbJMNqPQmX8vmLh0v/9BEd
AA4BAn1tFVEwoHh81olO97kvIxMCyEIHEzOwgLwYhR/3ifNu6cFH7N6+PeQikvM78srlzhcoHD7f
XUzEhugJzlVSb7ZPR3puiAsjRJ8yA7tbuJStOfRUpQ+yhBnVyXMpiaQ2Rb+aYiSRQOTdDYc7JcTG
GM4+HIuu6kgtI5IZwkdgJnawfJRz8BA3GM9JfdpWlxoSb8MS+DcAAcAdlAT7iIQEJAAwWFOKmqA4
IDgECYs1Vx0e3fGbLQXnvQLE6YZcmmdc7vkHXMCIZb0vGKaJUJWmEClJVSG7vAKQiBFENdsyn/Az
sWAT+JM/bCKp4Aw7aAv5WomSY0vcj+M3qaF4oXnf19dx9r6bwfWO8sY8RxgoE0Jqzl6KEUHq2pFq
UFuytGL/l2xGQRi3CL+PzXh6OdINPwof7iSIz56bhfYz+gX1RKzYGRhVb5gNH/eDyHM1FWwC14xH
/urtJUMZ5WMKe7XnO7B69vk5qBMTcZD2NdZD/uJBrWL4sNyFhUtnueijNRUwUPJN8vw7dF3/+wpr
6x/a+cG6Oyy6wolHbg0DZ8d6e6DLO6egNZxsNcTHylgiWx23SnGpBmmV5oRJuOY8Ekvr4JczRVPx
4A7nuGiu2ihkFFX+AG8szfMu65Glr2XOU2XFk9fYqrH6gOVg
`protect end_protected
